MACRO tl_synth_v4
  CLASS BLOCK ;
  FOREIGN tl_synth_v4 ;
  ORIGIN -284.500 -104.000 ;
  SIZE 142.500 BY 196.000 ;
  PIN VDD
    ANTENNAGATEAREA 66.423500 ;
    ANTENNADIFFAREA 179.243042 ;
    PORT
      LAYER met1 ;
        RECT 284.500 200.000 288.500 204.000 ;
    END
  END VDD
  PIN VSS
    ANTENNAGATEAREA 105.069901 ;
    ANTENNADIFFAREA 440.560547 ;
    PORT
      LAYER met1 ;
        RECT 284.500 205.000 288.500 209.000 ;
    END
  END VSS
  PIN VFREF
    ANTENNAGATEAREA 3.600000 ;
    PORT
      LAYER met3 ;
        RECT 284.500 190.250 286.500 192.250 ;
    END
  END VFREF
  PIN DI_DIV_N_CON[3]
    ANTENNAGATEAREA 0.607500 ;
    PORT
      LAYER met3 ;
        RECT 284.500 149.500 285.500 150.500 ;
    END
  END DI_DIV_N_CON[3]
  PIN DI_DIV_N_CON[2]
    ANTENNAGATEAREA 0.607500 ;
    PORT
      LAYER met3 ;
        RECT 284.500 148.000 285.500 149.000 ;
    END
  END DI_DIV_N_CON[2]
  PIN DI_DIV_N_CON[1]
    ANTENNAGATEAREA 0.607500 ;
    PORT
      LAYER met3 ;
        RECT 284.500 146.500 285.500 147.500 ;
    END
  END DI_DIV_N_CON[1]
  PIN DI_DIV_N_CON[0]
    ANTENNAGATEAREA 0.607500 ;
    PORT
      LAYER met3 ;
        RECT 284.500 145.000 285.500 146.000 ;
    END
  END DI_DIV_N_CON[0]
  PIN VCON_VCO
    ANTENNADIFFAREA 40.340000 ;
    PORT
      LAYER met3 ;
        RECT 376.000 157.500 377.500 159.000 ;
    END
  END VCON_VCO
  PIN DI_VCO_DISCRETE_CON[0]
    ANTENNAGATEAREA 1.737000 ;
    PORT
      LAYER met3 ;
        RECT 284.500 182.500 285.500 183.500 ;
    END
  END DI_VCO_DISCRETE_CON[0]
  PIN DI_VCO_DISCRETE_CON[1]
    ANTENNAGATEAREA 1.737000 ;
    PORT
      LAYER met3 ;
        RECT 284.500 181.000 285.500 182.000 ;
    END
  END DI_VCO_DISCRETE_CON[1]
  PIN DI_VCO_DISCRETE_CON[2]
    ANTENNAGATEAREA 1.494000 ;
    PORT
      LAYER met3 ;
        RECT 284.500 179.500 285.500 180.500 ;
    END
  END DI_VCO_DISCRETE_CON[2]
  PIN DI_VCO_DISCRETE_CON[3]
    ANTENNAGATEAREA 1.900500 ;
    PORT
      LAYER met3 ;
        RECT 284.500 178.000 285.500 179.000 ;
    END
  END DI_VCO_DISCRETE_CON[3]
  PIN VFOUT_HF
    ANTENNADIFFAREA 0.391500 ;
    PORT
      LAYER met3 ;
        RECT 284.500 117.750 285.500 118.750 ;
    END
  END VFOUT_HF
  PIN VFOUT_LF
    ANTENNADIFFAREA 0.391500 ;
    PORT
      LAYER met3 ;
        RECT 284.500 119.750 285.500 120.750 ;
    END
  END VFOUT_LF
  OBS
      LAYER nwell ;
        RECT 325.695 192.445 343.805 198.305 ;
      LAYER pwell ;
        RECT 325.695 184.195 343.805 189.305 ;
        RECT 349.000 189.000 356.000 193.500 ;
      LAYER nwell ;
        RECT 292.830 181.945 317.590 183.550 ;
      LAYER pwell ;
        RECT 293.025 180.745 294.395 181.555 ;
        RECT 294.405 180.745 299.915 181.555 ;
        RECT 299.925 180.745 305.435 181.555 ;
        RECT 305.915 180.830 306.345 181.615 ;
        RECT 306.365 180.745 311.875 181.555 ;
        RECT 311.885 180.745 315.555 181.555 ;
        RECT 316.025 180.745 317.395 181.555 ;
        RECT 293.165 180.535 293.335 180.745 ;
        RECT 294.545 180.535 294.715 180.745 ;
        RECT 297.300 180.585 297.420 180.695 ;
        RECT 300.065 180.555 300.235 180.745 ;
        RECT 300.065 180.535 300.205 180.555 ;
        RECT 300.525 180.535 300.695 180.725 ;
        RECT 305.580 180.585 305.700 180.695 ;
        RECT 306.045 180.535 306.215 180.725 ;
        RECT 306.505 180.555 306.675 180.745 ;
        RECT 312.025 180.555 312.195 180.745 ;
        RECT 314.320 180.535 314.490 180.725 ;
        RECT 314.785 180.535 314.955 180.725 ;
        RECT 315.700 180.585 315.820 180.695 ;
        RECT 317.085 180.535 317.255 180.745 ;
        RECT 293.025 179.725 294.395 180.535 ;
        RECT 294.405 179.725 297.155 180.535 ;
        RECT 297.635 179.715 300.205 180.535 ;
        RECT 300.385 179.725 305.895 180.535 ;
        RECT 305.905 179.725 311.415 180.535 ;
        RECT 297.635 179.625 299.225 179.715 ;
        RECT 311.425 179.625 314.635 180.535 ;
        RECT 314.645 179.725 316.015 180.535 ;
        RECT 316.025 179.725 317.395 180.535 ;
      LAYER nwell ;
        RECT 292.830 176.505 317.590 179.335 ;
      LAYER pwell ;
        RECT 293.025 175.305 294.395 176.115 ;
        RECT 294.405 175.305 295.775 176.115 ;
        RECT 295.785 175.305 298.995 176.215 ;
        RECT 299.910 175.985 301.280 176.215 ;
        RECT 299.005 175.305 301.280 175.985 ;
        RECT 301.305 175.305 304.975 176.115 ;
        RECT 305.915 175.390 306.345 176.175 ;
        RECT 306.365 175.305 310.035 176.115 ;
        RECT 310.965 175.305 314.175 176.215 ;
        RECT 314.185 175.305 316.015 176.115 ;
        RECT 316.025 175.305 317.395 176.115 ;
        RECT 293.165 175.095 293.335 175.305 ;
        RECT 294.545 175.095 294.715 175.305 ;
        RECT 295.930 175.285 296.100 175.305 ;
        RECT 295.925 175.115 296.100 175.285 ;
        RECT 293.025 174.285 294.395 175.095 ;
        RECT 294.405 174.285 295.775 175.095 ;
        RECT 295.925 175.065 296.095 175.115 ;
        RECT 298.685 175.095 298.855 175.285 ;
        RECT 299.150 175.115 299.320 175.305 ;
        RECT 301.445 175.115 301.615 175.305 ;
        RECT 304.205 175.095 304.375 175.285 ;
        RECT 305.135 175.150 305.295 175.260 ;
        RECT 306.505 175.115 306.675 175.305 ;
        RECT 309.725 175.095 309.895 175.285 ;
        RECT 310.195 175.150 310.355 175.260 ;
        RECT 313.860 175.115 314.030 175.305 ;
        RECT 314.325 175.115 314.495 175.305 ;
        RECT 315.255 175.140 315.415 175.250 ;
        RECT 317.085 175.095 317.255 175.305 ;
        RECT 297.125 175.065 298.505 175.095 ;
        RECT 295.800 174.385 298.505 175.065 ;
        RECT 297.125 174.185 298.505 174.385 ;
        RECT 298.545 174.285 304.055 175.095 ;
        RECT 304.065 174.285 309.575 175.095 ;
        RECT 309.585 174.285 315.095 175.095 ;
        RECT 316.025 174.285 317.395 175.095 ;
      LAYER nwell ;
        RECT 292.830 171.065 317.590 173.895 ;
      LAYER pwell ;
        RECT 293.025 169.865 294.395 170.675 ;
        RECT 294.405 169.865 296.235 170.675 ;
        RECT 296.705 169.865 299.915 170.775 ;
        RECT 299.925 169.865 305.435 170.675 ;
        RECT 305.915 169.950 306.345 170.735 ;
        RECT 306.365 169.865 310.035 170.675 ;
        RECT 310.045 169.865 311.415 170.675 ;
        RECT 311.425 169.865 314.465 170.775 ;
        RECT 314.645 169.865 316.015 170.675 ;
        RECT 316.025 169.865 317.395 170.675 ;
        RECT 293.165 169.655 293.335 169.865 ;
        RECT 294.545 169.655 294.715 169.865 ;
        RECT 296.380 169.705 296.500 169.815 ;
        RECT 296.850 169.675 297.020 169.865 ;
        RECT 300.065 169.655 300.235 169.865 ;
        RECT 305.585 169.815 305.755 169.845 ;
        RECT 305.580 169.705 305.755 169.815 ;
        RECT 305.585 169.655 305.755 169.705 ;
        RECT 306.505 169.675 306.675 169.865 ;
        RECT 310.185 169.675 310.355 169.865 ;
        RECT 314.320 169.845 314.465 169.865 ;
        RECT 311.105 169.655 311.275 169.845 ;
        RECT 312.485 169.655 312.655 169.845 ;
        RECT 314.320 169.675 314.495 169.845 ;
        RECT 314.785 169.675 314.955 169.865 ;
        RECT 314.325 169.655 314.495 169.675 ;
        RECT 317.085 169.655 317.255 169.865 ;
        RECT 293.025 168.845 294.395 169.655 ;
        RECT 294.405 168.845 299.915 169.655 ;
        RECT 299.925 168.845 305.435 169.655 ;
        RECT 305.445 168.845 310.955 169.655 ;
        RECT 310.965 168.845 312.335 169.655 ;
        RECT 312.345 168.975 314.175 169.655 ;
        RECT 312.830 168.745 314.175 168.975 ;
        RECT 314.185 168.845 316.015 169.655 ;
        RECT 316.025 168.845 317.395 169.655 ;
      LAYER nwell ;
        RECT 292.830 165.625 317.590 168.455 ;
      LAYER pwell ;
        RECT 387.750 166.000 391.750 197.000 ;
        RECT 397.250 166.000 401.250 197.000 ;
        RECT 406.750 166.000 410.750 197.000 ;
        RECT 293.025 164.425 294.395 165.235 ;
        RECT 294.405 164.425 297.155 165.235 ;
        RECT 297.640 165.105 299.010 165.335 ;
        RECT 300.385 165.135 301.795 165.335 ;
        RECT 297.640 164.425 299.915 165.105 ;
        RECT 300.385 164.455 303.120 165.135 ;
        RECT 300.385 164.425 301.780 164.455 ;
        RECT 293.165 164.215 293.335 164.425 ;
        RECT 294.545 164.235 294.715 164.425 ;
        RECT 295.465 164.235 295.635 164.405 ;
        RECT 295.930 164.235 296.100 164.405 ;
        RECT 297.300 164.265 297.420 164.375 ;
        RECT 299.600 164.235 299.770 164.425 ;
        RECT 300.060 164.265 300.180 164.375 ;
        RECT 301.445 164.235 301.615 164.405 ;
        RECT 295.955 164.215 296.100 164.235 ;
        RECT 301.445 164.215 301.585 164.235 ;
        RECT 301.905 164.215 302.075 164.405 ;
        RECT 302.825 164.235 302.995 164.455 ;
        RECT 303.145 164.425 305.895 165.235 ;
        RECT 305.915 164.510 306.345 165.295 ;
        RECT 306.365 164.425 310.035 165.235 ;
        RECT 310.505 164.425 313.545 165.335 ;
        RECT 313.725 164.425 315.555 165.235 ;
        RECT 316.025 164.425 317.395 165.235 ;
        RECT 303.285 164.235 303.455 164.425 ;
        RECT 306.505 164.235 306.675 164.425 ;
        RECT 313.400 164.405 313.545 164.425 ;
        RECT 307.425 164.215 307.595 164.405 ;
        RECT 310.180 164.265 310.300 164.375 ;
        RECT 311.100 164.265 311.220 164.375 ;
        RECT 313.400 164.235 313.570 164.405 ;
        RECT 313.865 164.235 314.035 164.425 ;
        RECT 314.320 164.235 314.490 164.405 ;
        RECT 314.320 164.215 314.465 164.235 ;
        RECT 314.785 164.215 314.955 164.405 ;
        RECT 315.700 164.265 315.820 164.375 ;
        RECT 317.085 164.215 317.255 164.425 ;
        RECT 293.025 163.405 294.395 164.215 ;
        RECT 295.955 163.305 298.995 164.215 ;
        RECT 299.015 163.395 301.585 164.215 ;
        RECT 301.765 163.405 307.275 164.215 ;
        RECT 307.285 163.405 310.955 164.215 ;
        RECT 299.015 163.305 300.605 163.395 ;
        RECT 311.425 163.305 314.465 164.215 ;
        RECT 314.645 163.405 316.015 164.215 ;
        RECT 316.025 163.405 317.395 164.215 ;
      LAYER nwell ;
        RECT 292.830 160.185 317.590 163.015 ;
      LAYER pwell ;
        RECT 293.025 158.985 294.395 159.795 ;
        RECT 294.405 158.985 299.915 159.795 ;
        RECT 299.925 158.985 305.435 159.795 ;
        RECT 305.915 159.070 306.345 159.855 ;
        RECT 306.365 158.985 311.875 159.795 ;
        RECT 311.885 158.985 315.555 159.795 ;
        RECT 316.025 158.985 317.395 159.795 ;
        RECT 293.165 158.795 293.335 158.985 ;
        RECT 294.545 158.795 294.715 158.985 ;
        RECT 300.065 158.795 300.235 158.985 ;
        RECT 305.580 158.825 305.700 158.935 ;
        RECT 306.505 158.795 306.675 158.985 ;
        RECT 312.025 158.795 312.195 158.985 ;
        RECT 315.700 158.825 315.820 158.935 ;
        RECT 317.085 158.795 317.255 158.985 ;
        RECT 379.000 158.250 390.500 164.250 ;
      LAYER nwell ;
        RECT 390.500 163.750 409.500 165.750 ;
        RECT 390.500 158.250 421.250 163.750 ;
      LAYER pwell ;
        RECT 379.000 152.750 421.250 158.250 ;
        RECT 379.000 152.250 409.500 152.750 ;
        RECT 390.500 150.750 409.500 152.250 ;
      LAYER nwell ;
        RECT 287.250 146.185 344.500 147.705 ;
      LAYER pwell ;
        RECT 287.250 145.770 344.500 145.855 ;
        RECT 287.250 145.730 287.430 145.770 ;
        RECT 287.750 145.730 301.430 145.770 ;
        RECT 301.820 145.730 313.930 145.770 ;
        RECT 314.320 145.730 323.930 145.770 ;
        RECT 324.320 145.730 334.680 145.770 ;
        RECT 335.070 145.730 343.930 145.770 ;
        RECT 344.320 145.730 344.500 145.770 ;
        RECT 287.250 144.785 344.500 145.730 ;
      LAYER nwell ;
        RECT 293.000 139.185 341.250 140.705 ;
        RECT 343.500 139.185 351.000 140.705 ;
      LAYER pwell ;
        RECT 293.000 138.770 341.250 138.855 ;
        RECT 293.000 138.730 293.180 138.770 ;
        RECT 293.570 138.730 298.180 138.770 ;
        RECT 298.570 138.730 303.180 138.770 ;
        RECT 303.570 138.730 310.930 138.770 ;
        RECT 311.320 138.730 320.680 138.770 ;
        RECT 321.070 138.730 327.680 138.770 ;
        RECT 328.070 138.730 333.680 138.770 ;
        RECT 334.070 138.730 340.680 138.770 ;
        RECT 341.070 138.730 341.250 138.770 ;
        RECT 293.000 137.785 341.250 138.730 ;
        RECT 343.500 138.770 351.000 138.855 ;
        RECT 343.500 138.730 348.680 138.770 ;
        RECT 349.070 138.730 351.000 138.770 ;
        RECT 343.500 137.785 351.000 138.730 ;
      LAYER nwell ;
        RECT 292.750 132.185 351.000 133.705 ;
      LAYER pwell ;
        RECT 292.750 131.770 351.000 131.855 ;
        RECT 292.750 131.730 292.930 131.770 ;
        RECT 293.320 131.730 303.180 131.770 ;
        RECT 303.570 131.730 310.930 131.770 ;
        RECT 311.320 131.730 315.430 131.770 ;
        RECT 315.820 131.730 322.430 131.770 ;
        RECT 322.820 131.730 328.430 131.770 ;
        RECT 328.820 131.730 335.430 131.770 ;
        RECT 335.820 131.730 341.430 131.770 ;
        RECT 341.820 131.730 348.680 131.770 ;
        RECT 349.070 131.730 351.000 131.770 ;
        RECT 292.750 130.785 351.000 131.730 ;
      LAYER nwell ;
        RECT 298.500 121.935 346.500 123.455 ;
      LAYER pwell ;
        RECT 298.500 121.520 346.500 121.605 ;
        RECT 298.500 121.480 307.180 121.520 ;
        RECT 307.570 121.480 323.180 121.520 ;
        RECT 323.570 121.480 339.180 121.520 ;
        RECT 339.570 121.480 346.500 121.520 ;
        RECT 298.500 120.535 346.500 121.480 ;
        RECT 387.750 119.500 391.750 150.500 ;
        RECT 397.250 119.500 401.250 150.500 ;
        RECT 406.750 119.500 410.750 150.500 ;
      LAYER nwell ;
        RECT 298.500 115.685 346.000 117.205 ;
      LAYER pwell ;
        RECT 298.500 115.270 346.000 115.355 ;
        RECT 298.500 115.230 300.430 115.270 ;
        RECT 300.820 115.230 306.180 115.270 ;
        RECT 306.570 115.230 306.930 115.270 ;
        RECT 307.320 115.230 307.680 115.270 ;
        RECT 308.000 115.230 313.180 115.270 ;
        RECT 313.570 115.230 313.930 115.270 ;
        RECT 314.320 115.230 316.430 115.270 ;
        RECT 316.820 115.230 326.930 115.270 ;
        RECT 327.320 115.230 332.430 115.270 ;
        RECT 332.820 115.230 338.180 115.270 ;
        RECT 338.570 115.230 338.930 115.270 ;
        RECT 339.320 115.230 344.680 115.270 ;
        RECT 345.070 115.230 345.430 115.270 ;
        RECT 345.820 115.230 346.000 115.270 ;
        RECT 298.500 114.285 346.000 115.230 ;
      LAYER li1 ;
        RECT 325.875 197.875 343.625 198.125 ;
        RECT 325.875 192.875 326.125 197.875 ;
        RECT 326.555 194.620 326.725 196.660 ;
        RECT 326.995 194.620 327.165 196.660 ;
        RECT 327.435 194.620 327.605 196.660 ;
        RECT 327.875 194.620 328.045 196.660 ;
        RECT 328.315 194.620 328.485 196.660 ;
        RECT 328.965 194.620 329.135 196.660 ;
        RECT 329.405 194.620 329.575 196.660 ;
        RECT 329.845 194.620 330.015 196.660 ;
        RECT 330.285 194.620 330.455 196.660 ;
        RECT 330.725 194.620 330.895 196.660 ;
        RECT 331.375 194.620 331.545 196.660 ;
        RECT 331.815 194.620 331.985 196.660 ;
        RECT 332.255 194.620 332.425 196.660 ;
        RECT 332.695 194.620 332.865 196.660 ;
        RECT 333.135 194.620 333.305 196.660 ;
        RECT 333.785 194.620 333.955 196.660 ;
        RECT 334.225 194.620 334.395 196.660 ;
        RECT 334.665 194.620 334.835 196.660 ;
        RECT 335.105 194.620 335.275 196.660 ;
        RECT 335.545 194.620 335.715 196.660 ;
        RECT 336.195 194.620 336.365 196.660 ;
        RECT 336.635 194.620 336.805 196.660 ;
        RECT 337.075 194.620 337.245 196.660 ;
        RECT 337.515 194.620 337.685 196.660 ;
        RECT 337.955 194.620 338.125 196.660 ;
        RECT 338.605 194.620 338.775 196.660 ;
        RECT 339.045 194.620 339.215 196.660 ;
        RECT 339.485 194.620 339.655 196.660 ;
        RECT 339.925 194.620 340.095 196.660 ;
        RECT 340.365 194.620 340.535 196.660 ;
        RECT 341.015 194.620 341.185 196.660 ;
        RECT 341.455 194.620 341.625 196.660 ;
        RECT 341.895 194.620 342.065 196.660 ;
        RECT 342.335 194.620 342.505 196.660 ;
        RECT 342.775 194.620 342.945 196.660 ;
        RECT 327.355 193.310 327.685 193.690 ;
        RECT 329.765 193.310 330.095 193.690 ;
        RECT 332.175 193.310 332.505 193.690 ;
        RECT 334.585 193.310 334.915 193.690 ;
        RECT 336.995 193.310 337.325 193.690 ;
        RECT 339.405 193.310 339.735 193.690 ;
        RECT 341.815 193.310 342.145 193.690 ;
        RECT 343.375 192.875 343.625 197.875 ;
        RECT 388.125 196.375 391.375 196.625 ;
        RECT 325.875 192.625 343.625 192.875 ;
        RECT 349.375 192.875 355.625 193.125 ;
        RECT 349.375 189.625 349.625 192.875 ;
        RECT 350.835 192.030 351.165 192.470 ;
        RECT 350.425 190.730 350.865 191.770 ;
        RECT 351.135 190.730 351.575 191.770 ;
        RECT 350.835 190.030 351.165 190.470 ;
        RECT 352.375 189.625 352.625 192.875 ;
        RECT 353.835 192.030 354.165 192.470 ;
        RECT 353.425 190.730 353.865 191.770 ;
        RECT 354.135 190.730 354.575 191.770 ;
        RECT 353.835 190.030 354.165 190.470 ;
        RECT 355.375 189.625 355.625 192.875 ;
        RECT 349.375 189.375 355.625 189.625 ;
        RECT 388.125 192.875 388.375 196.375 ;
        RECT 389.665 195.250 389.835 195.750 ;
        RECT 388.780 193.980 389.260 195.020 ;
        RECT 389.530 193.980 389.970 195.020 ;
        RECT 390.240 193.980 390.720 195.020 ;
        RECT 389.665 193.250 389.835 193.750 ;
        RECT 391.125 192.875 391.375 196.375 ;
        RECT 388.125 192.625 391.375 192.875 ;
        RECT 388.125 189.125 388.375 192.625 ;
        RECT 389.665 191.500 389.835 192.000 ;
        RECT 388.780 190.230 389.260 191.270 ;
        RECT 389.530 190.230 389.970 191.270 ;
        RECT 390.240 190.230 390.720 191.270 ;
        RECT 389.665 189.500 389.835 190.000 ;
        RECT 391.125 189.125 391.375 192.625 ;
        RECT 325.875 188.875 343.625 189.125 ;
        RECT 325.875 184.625 326.125 188.875 ;
        RECT 327.355 188.060 327.685 188.440 ;
        RECT 329.765 188.060 330.095 188.440 ;
        RECT 332.175 188.060 332.505 188.440 ;
        RECT 334.585 188.060 334.915 188.440 ;
        RECT 336.995 188.060 337.325 188.440 ;
        RECT 339.405 188.060 339.735 188.440 ;
        RECT 341.815 188.060 342.145 188.440 ;
        RECT 326.555 186.090 326.725 187.130 ;
        RECT 326.995 186.090 327.165 187.130 ;
        RECT 327.435 186.090 327.605 187.130 ;
        RECT 327.875 186.090 328.045 187.130 ;
        RECT 328.315 186.090 328.485 187.130 ;
        RECT 328.965 186.090 329.135 187.130 ;
        RECT 329.405 186.090 329.575 187.130 ;
        RECT 329.845 186.090 330.015 187.130 ;
        RECT 330.285 186.090 330.455 187.130 ;
        RECT 330.725 186.090 330.895 187.130 ;
        RECT 331.375 186.090 331.545 187.130 ;
        RECT 331.815 186.090 331.985 187.130 ;
        RECT 332.255 186.090 332.425 187.130 ;
        RECT 332.695 186.090 332.865 187.130 ;
        RECT 333.135 186.090 333.305 187.130 ;
        RECT 333.785 186.090 333.955 187.130 ;
        RECT 334.225 186.090 334.395 187.130 ;
        RECT 334.665 186.090 334.835 187.130 ;
        RECT 335.105 186.090 335.275 187.130 ;
        RECT 335.545 186.090 335.715 187.130 ;
        RECT 336.195 186.090 336.365 187.130 ;
        RECT 336.635 186.090 336.805 187.130 ;
        RECT 337.075 186.090 337.245 187.130 ;
        RECT 337.515 186.090 337.685 187.130 ;
        RECT 337.955 186.090 338.125 187.130 ;
        RECT 338.605 186.090 338.775 187.130 ;
        RECT 339.045 186.090 339.215 187.130 ;
        RECT 339.485 186.090 339.655 187.130 ;
        RECT 339.925 186.090 340.095 187.130 ;
        RECT 340.365 186.090 340.535 187.130 ;
        RECT 341.015 186.090 341.185 187.130 ;
        RECT 341.455 186.090 341.625 187.130 ;
        RECT 341.895 186.090 342.065 187.130 ;
        RECT 342.335 186.090 342.505 187.130 ;
        RECT 342.775 186.090 342.945 187.130 ;
        RECT 343.375 184.625 343.625 188.875 ;
        RECT 325.875 184.375 343.625 184.625 ;
        RECT 388.125 188.875 391.375 189.125 ;
        RECT 388.125 185.375 388.375 188.875 ;
        RECT 389.665 187.750 389.835 188.250 ;
        RECT 388.780 186.480 389.260 187.520 ;
        RECT 389.530 186.480 389.970 187.520 ;
        RECT 390.240 186.480 390.720 187.520 ;
        RECT 389.665 185.750 389.835 186.250 ;
        RECT 391.125 185.375 391.375 188.875 ;
        RECT 388.125 185.125 391.375 185.375 ;
        RECT 293.020 183.275 317.400 183.445 ;
        RECT 293.105 182.185 294.315 183.275 ;
        RECT 294.485 182.840 299.830 183.275 ;
        RECT 300.005 182.840 305.350 183.275 ;
        RECT 293.105 181.475 293.625 182.015 ;
        RECT 293.795 181.645 294.315 182.185 ;
        RECT 293.105 180.725 294.315 181.475 ;
        RECT 296.070 181.270 296.410 182.100 ;
        RECT 297.890 181.590 298.240 182.840 ;
        RECT 301.590 181.270 301.930 182.100 ;
        RECT 303.410 181.590 303.760 182.840 ;
        RECT 305.985 182.110 306.275 183.275 ;
        RECT 306.445 182.840 311.790 183.275 ;
        RECT 294.485 180.725 299.830 181.270 ;
        RECT 300.005 180.725 305.350 181.270 ;
        RECT 305.985 180.725 306.275 181.450 ;
        RECT 308.030 181.270 308.370 182.100 ;
        RECT 309.850 181.590 310.200 182.840 ;
        RECT 311.965 182.185 315.475 183.275 ;
        RECT 311.965 181.495 313.615 182.015 ;
        RECT 313.785 181.665 315.475 182.185 ;
        RECT 316.105 182.185 317.315 183.275 ;
        RECT 316.105 181.645 316.625 182.185 ;
        RECT 306.445 180.725 311.790 181.270 ;
        RECT 311.965 180.725 315.475 181.495 ;
        RECT 316.795 181.475 317.315 182.015 ;
        RECT 316.105 180.725 317.315 181.475 ;
        RECT 388.125 181.625 388.375 185.125 ;
        RECT 389.665 184.000 389.835 184.500 ;
        RECT 388.780 182.730 389.260 183.770 ;
        RECT 389.530 182.730 389.970 183.770 ;
        RECT 390.240 182.730 390.720 183.770 ;
        RECT 389.665 182.000 389.835 182.500 ;
        RECT 391.125 181.625 391.375 185.125 ;
        RECT 388.125 181.375 391.375 181.625 ;
        RECT 293.020 180.555 317.400 180.725 ;
        RECT 293.105 179.805 294.315 180.555 ;
        RECT 293.105 179.265 293.625 179.805 ;
        RECT 294.485 179.785 297.075 180.555 ;
        RECT 293.795 179.095 294.315 179.635 ;
        RECT 294.485 179.265 295.695 179.785 ;
        RECT 297.705 179.755 297.995 180.555 ;
        RECT 298.165 180.095 298.715 180.385 ;
        RECT 298.885 180.095 299.135 180.555 ;
        RECT 295.865 179.095 297.075 179.615 ;
        RECT 293.105 178.005 294.315 179.095 ;
        RECT 294.485 178.005 297.075 179.095 ;
        RECT 297.705 178.005 297.995 179.145 ;
        RECT 298.165 178.725 298.415 180.095 ;
        RECT 299.765 179.925 300.095 180.285 ;
        RECT 300.465 180.010 305.810 180.555 ;
        RECT 305.985 180.010 311.330 180.555 ;
        RECT 311.505 180.075 311.765 180.555 ;
        RECT 311.935 180.305 312.180 180.385 ;
        RECT 311.935 180.135 312.265 180.305 ;
        RECT 298.705 179.735 300.095 179.925 ;
        RECT 298.705 179.645 298.875 179.735 ;
        RECT 298.585 179.315 298.875 179.645 ;
        RECT 299.045 179.315 299.375 179.565 ;
        RECT 299.605 179.315 300.295 179.565 ;
        RECT 298.705 179.065 298.875 179.315 ;
        RECT 298.705 178.895 299.645 179.065 ;
        RECT 298.165 178.175 298.615 178.725 ;
        RECT 298.805 178.005 299.135 178.725 ;
        RECT 299.345 178.345 299.645 178.895 ;
        RECT 299.980 178.875 300.295 179.315 ;
        RECT 302.050 179.180 302.390 180.010 ;
        RECT 299.815 178.005 300.095 178.675 ;
        RECT 303.870 178.440 304.220 179.690 ;
        RECT 307.570 179.180 307.910 180.010 ;
        RECT 309.390 178.440 309.740 179.690 ;
        RECT 311.550 179.315 311.745 179.885 ;
        RECT 311.935 179.145 312.105 180.135 ;
        RECT 312.465 179.940 312.675 180.225 ;
        RECT 312.940 180.215 313.110 180.240 ;
        RECT 312.940 180.045 313.115 180.215 ;
        RECT 313.355 180.175 313.685 180.555 ;
        RECT 313.455 180.095 313.625 180.175 ;
        RECT 312.940 179.945 313.110 180.045 ;
        RECT 312.285 179.770 312.675 179.940 ;
        RECT 312.845 179.775 313.110 179.945 ;
        RECT 313.875 179.925 314.045 180.385 ;
        RECT 314.295 180.095 314.550 180.555 ;
        RECT 312.285 179.315 312.455 179.770 ;
        RECT 312.845 179.565 313.015 179.775 ;
        RECT 313.370 179.645 313.575 179.880 ;
        RECT 313.875 179.755 314.550 179.925 ;
        RECT 312.685 179.395 313.015 179.565 ;
        RECT 312.845 179.380 313.015 179.395 ;
        RECT 313.245 179.315 313.575 179.645 ;
        RECT 313.755 179.395 314.085 179.565 ;
        RECT 313.915 179.145 314.085 179.395 ;
        RECT 311.595 178.975 314.085 179.145 ;
        RECT 300.465 178.005 305.810 178.440 ;
        RECT 305.985 178.005 311.330 178.440 ;
        RECT 311.595 178.175 311.765 178.975 ;
        RECT 314.295 178.805 314.550 179.755 ;
        RECT 314.725 179.805 315.935 180.555 ;
        RECT 316.105 179.805 317.315 180.555 ;
        RECT 314.725 179.265 315.245 179.805 ;
        RECT 315.415 179.095 315.935 179.635 ;
        RECT 311.995 178.635 313.285 178.805 ;
        RECT 312.055 178.215 312.305 178.635 ;
        RECT 312.495 178.005 312.825 178.465 ;
        RECT 313.035 178.215 313.285 178.635 ;
        RECT 313.455 178.005 313.705 178.805 ;
        RECT 313.875 178.635 314.550 178.805 ;
        RECT 313.875 178.175 314.045 178.635 ;
        RECT 314.255 178.005 314.505 178.465 ;
        RECT 314.725 178.005 315.935 179.095 ;
        RECT 316.105 179.095 316.625 179.635 ;
        RECT 316.795 179.265 317.315 179.805 ;
        RECT 316.105 178.005 317.315 179.095 ;
        RECT 293.020 177.835 317.400 178.005 ;
        RECT 388.125 177.875 388.375 181.375 ;
        RECT 389.665 180.250 389.835 180.750 ;
        RECT 388.780 178.980 389.260 180.020 ;
        RECT 389.530 178.980 389.970 180.020 ;
        RECT 390.240 178.980 390.720 180.020 ;
        RECT 389.665 178.250 389.835 178.750 ;
        RECT 391.125 177.875 391.375 181.375 ;
        RECT 293.105 176.745 294.315 177.835 ;
        RECT 294.485 176.745 295.695 177.835 ;
        RECT 295.915 177.375 296.165 177.835 ;
        RECT 296.375 177.205 296.545 177.665 ;
        RECT 293.105 176.035 293.625 176.575 ;
        RECT 293.795 176.205 294.315 176.745 ;
        RECT 294.485 176.035 295.005 176.575 ;
        RECT 295.175 176.205 295.695 176.745 ;
        RECT 295.870 177.035 296.545 177.205 ;
        RECT 296.715 177.035 296.965 177.835 ;
        RECT 297.135 177.205 297.385 177.625 ;
        RECT 297.595 177.375 297.925 177.835 ;
        RECT 298.115 177.205 298.365 177.625 ;
        RECT 297.135 177.035 298.425 177.205 ;
        RECT 295.870 176.085 296.125 177.035 ;
        RECT 298.655 176.865 298.825 177.665 ;
        RECT 296.335 176.695 298.825 176.865 ;
        RECT 299.155 176.865 299.515 177.040 ;
        RECT 300.100 177.035 300.270 177.835 ;
        RECT 300.440 177.205 300.770 177.665 ;
        RECT 300.940 177.375 301.110 177.835 ;
        RECT 300.440 177.035 301.215 177.205 ;
        RECT 299.155 176.695 300.615 176.865 ;
        RECT 296.335 176.445 296.505 176.695 ;
        RECT 296.335 176.275 296.665 176.445 ;
        RECT 296.845 176.195 297.175 176.525 ;
        RECT 297.405 176.445 297.575 176.460 ;
        RECT 297.405 176.275 297.735 176.445 ;
        RECT 293.105 175.285 294.315 176.035 ;
        RECT 294.485 175.285 295.695 176.035 ;
        RECT 295.870 175.915 296.545 176.085 ;
        RECT 296.845 175.960 297.050 176.195 ;
        RECT 297.405 176.065 297.575 176.275 ;
        RECT 297.965 176.070 298.135 176.525 ;
        RECT 295.870 175.285 296.125 175.745 ;
        RECT 296.375 175.455 296.545 175.915 ;
        RECT 297.310 175.895 297.575 176.065 ;
        RECT 297.745 175.900 298.135 176.070 ;
        RECT 297.310 175.795 297.480 175.895 ;
        RECT 296.795 175.665 296.965 175.745 ;
        RECT 296.735 175.285 297.065 175.665 ;
        RECT 297.305 175.625 297.480 175.795 ;
        RECT 297.310 175.600 297.480 175.625 ;
        RECT 297.745 175.615 297.955 175.900 ;
        RECT 298.315 175.705 298.485 176.695 ;
        RECT 298.675 175.955 298.870 176.525 ;
        RECT 299.150 176.475 299.345 176.525 ;
        RECT 299.145 176.305 299.345 176.475 ;
        RECT 299.150 175.965 299.345 176.305 ;
        RECT 299.515 175.795 299.695 176.695 ;
        RECT 299.865 175.965 300.275 176.525 ;
        RECT 300.445 176.195 300.615 176.695 ;
        RECT 300.785 176.025 301.215 177.035 ;
        RECT 301.385 176.745 304.895 177.835 ;
        RECT 300.520 175.855 301.215 176.025 ;
        RECT 301.385 176.055 303.035 176.575 ;
        RECT 303.205 176.225 304.895 176.745 ;
        RECT 305.985 176.670 306.275 177.835 ;
        RECT 306.445 176.745 309.955 177.835 ;
        RECT 311.060 176.850 311.385 177.835 ;
        RECT 311.955 177.205 312.215 177.665 ;
        RECT 312.385 177.385 313.235 177.835 ;
        RECT 311.570 177.155 311.775 177.185 ;
        RECT 311.565 176.985 311.775 177.155 ;
        RECT 311.955 176.985 313.075 177.205 ;
        RECT 306.445 176.055 308.095 176.575 ;
        RECT 308.265 176.225 309.955 176.745 ;
        RECT 311.055 176.195 311.315 176.650 ;
        RECT 311.570 176.600 311.775 176.985 ;
        RECT 311.570 176.225 312.155 176.600 ;
        RECT 312.325 176.210 312.735 176.815 ;
        RECT 312.905 176.530 313.075 176.985 ;
        RECT 298.155 175.535 298.485 175.705 ;
        RECT 298.240 175.455 298.485 175.535 ;
        RECT 298.655 175.285 298.915 175.765 ;
        RECT 299.105 175.285 299.345 175.795 ;
        RECT 299.515 175.455 299.805 175.795 ;
        RECT 300.035 175.285 300.350 175.795 ;
        RECT 300.520 175.585 300.690 175.855 ;
        RECT 300.860 175.285 301.190 175.685 ;
        RECT 301.385 175.285 304.895 176.055 ;
        RECT 305.985 175.285 306.275 176.010 ;
        RECT 306.445 175.285 309.955 176.055 ;
        RECT 312.905 176.040 313.235 176.530 ;
        RECT 311.060 175.835 312.215 176.025 ;
        RECT 311.060 175.695 311.335 175.835 ;
        RECT 312.005 175.665 312.215 175.835 ;
        RECT 312.385 175.835 313.235 176.040 ;
        RECT 311.505 175.285 311.835 175.665 ;
        RECT 312.385 175.455 312.715 175.835 ;
        RECT 312.905 175.285 313.235 175.665 ;
        RECT 313.405 175.455 313.650 177.665 ;
        RECT 313.835 176.835 314.090 177.835 ;
        RECT 314.265 176.745 315.935 177.835 ;
        RECT 313.835 175.285 314.075 176.085 ;
        RECT 314.265 176.055 315.015 176.575 ;
        RECT 315.185 176.225 315.935 176.745 ;
        RECT 316.105 176.745 317.315 177.835 ;
        RECT 388.125 177.625 391.375 177.875 ;
        RECT 316.105 176.205 316.625 176.745 ;
        RECT 314.265 175.285 315.935 176.055 ;
        RECT 316.795 176.035 317.315 176.575 ;
        RECT 316.105 175.285 317.315 176.035 ;
        RECT 293.020 175.115 317.400 175.285 ;
        RECT 293.105 174.365 294.315 175.115 ;
        RECT 294.485 174.365 295.695 175.115 ;
        RECT 295.885 174.545 296.140 174.895 ;
        RECT 296.310 174.715 296.640 175.115 ;
        RECT 296.810 174.545 296.980 174.895 ;
        RECT 297.150 174.715 297.530 175.115 ;
        RECT 295.885 174.375 297.550 174.545 ;
        RECT 297.720 174.440 297.995 174.785 ;
        RECT 293.105 173.825 293.625 174.365 ;
        RECT 293.795 173.655 294.315 174.195 ;
        RECT 294.485 173.825 295.005 174.365 ;
        RECT 297.380 174.205 297.550 174.375 ;
        RECT 295.175 173.655 295.695 174.195 ;
        RECT 295.865 173.875 296.215 174.205 ;
        RECT 296.385 173.875 297.210 174.205 ;
        RECT 297.380 173.875 297.655 174.205 ;
        RECT 293.105 172.565 294.315 173.655 ;
        RECT 294.485 172.565 295.695 173.655 ;
        RECT 295.885 173.415 296.215 173.705 ;
        RECT 296.385 173.585 296.610 173.875 ;
        RECT 297.380 173.705 297.550 173.875 ;
        RECT 297.825 173.705 297.995 174.440 ;
        RECT 298.165 174.285 298.455 175.115 ;
        RECT 298.625 174.570 303.970 175.115 ;
        RECT 304.145 174.570 309.490 175.115 ;
        RECT 309.665 174.570 315.010 175.115 ;
        RECT 296.880 173.535 297.550 173.705 ;
        RECT 296.880 173.415 297.050 173.535 ;
        RECT 295.885 173.245 297.050 173.415 ;
        RECT 295.865 172.785 297.060 173.075 ;
        RECT 297.230 172.565 297.510 173.365 ;
        RECT 297.720 172.735 297.995 173.705 ;
        RECT 298.165 172.565 298.455 173.770 ;
        RECT 300.210 173.740 300.550 174.570 ;
        RECT 302.030 173.000 302.380 174.250 ;
        RECT 305.730 173.740 306.070 174.570 ;
        RECT 307.550 173.000 307.900 174.250 ;
        RECT 311.250 173.740 311.590 174.570 ;
        RECT 316.105 174.365 317.315 175.115 ;
        RECT 313.070 173.000 313.420 174.250 ;
        RECT 316.105 173.655 316.625 174.195 ;
        RECT 316.795 173.825 317.315 174.365 ;
        RECT 388.125 174.125 388.375 177.625 ;
        RECT 389.665 176.500 389.835 177.000 ;
        RECT 388.780 175.230 389.260 176.270 ;
        RECT 389.530 175.230 389.970 176.270 ;
        RECT 390.240 175.230 390.720 176.270 ;
        RECT 389.665 174.500 389.835 175.000 ;
        RECT 391.125 174.125 391.375 177.625 ;
        RECT 388.125 173.875 391.375 174.125 ;
        RECT 298.625 172.565 303.970 173.000 ;
        RECT 304.145 172.565 309.490 173.000 ;
        RECT 309.665 172.565 315.010 173.000 ;
        RECT 316.105 172.565 317.315 173.655 ;
        RECT 293.020 172.395 317.400 172.565 ;
        RECT 293.105 171.305 294.315 172.395 ;
        RECT 294.485 171.305 296.155 172.395 ;
        RECT 296.790 171.395 297.045 172.395 ;
        RECT 293.105 170.595 293.625 171.135 ;
        RECT 293.795 170.765 294.315 171.305 ;
        RECT 294.485 170.615 295.235 171.135 ;
        RECT 295.405 170.785 296.155 171.305 ;
        RECT 293.105 169.845 294.315 170.595 ;
        RECT 294.485 169.845 296.155 170.615 ;
        RECT 296.805 169.845 297.045 170.645 ;
        RECT 297.230 170.015 297.475 172.225 ;
        RECT 297.645 171.945 298.495 172.395 ;
        RECT 298.665 171.765 298.925 172.225 ;
        RECT 297.805 171.545 298.925 171.765 ;
        RECT 299.105 171.715 299.310 171.745 ;
        RECT 299.105 171.545 299.315 171.715 ;
        RECT 297.805 171.090 297.975 171.545 ;
        RECT 297.645 170.600 297.975 171.090 ;
        RECT 298.145 170.770 298.555 171.375 ;
        RECT 299.105 171.160 299.310 171.545 ;
        RECT 299.495 171.410 299.820 172.395 ;
        RECT 300.005 171.960 305.350 172.395 ;
        RECT 298.725 170.785 299.310 171.160 ;
        RECT 299.565 170.755 299.825 171.210 ;
        RECT 297.645 170.395 298.495 170.600 ;
        RECT 297.645 169.845 297.975 170.225 ;
        RECT 298.165 170.015 298.495 170.395 ;
        RECT 298.665 170.395 299.820 170.585 ;
        RECT 298.665 170.225 298.875 170.395 ;
        RECT 299.545 170.255 299.820 170.395 ;
        RECT 301.590 170.390 301.930 171.220 ;
        RECT 303.410 170.710 303.760 171.960 ;
        RECT 305.985 171.230 306.275 172.395 ;
        RECT 306.445 171.305 309.955 172.395 ;
        RECT 310.125 171.305 311.335 172.395 ;
        RECT 311.565 171.695 311.785 172.225 ;
        RECT 311.955 171.885 312.285 172.395 ;
        RECT 312.455 171.695 312.680 172.225 ;
        RECT 311.565 171.430 312.680 171.695 ;
        RECT 312.850 171.680 313.165 172.225 ;
        RECT 313.355 171.980 313.685 172.395 ;
        RECT 312.850 171.450 313.685 171.680 ;
        RECT 306.445 170.615 308.095 171.135 ;
        RECT 308.265 170.785 309.955 171.305 ;
        RECT 299.045 169.845 299.375 170.225 ;
        RECT 300.005 169.845 305.350 170.390 ;
        RECT 305.985 169.845 306.275 170.570 ;
        RECT 306.445 169.845 309.955 170.615 ;
        RECT 310.125 170.595 310.645 171.135 ;
        RECT 310.815 170.765 311.335 171.305 ;
        RECT 310.125 169.845 311.335 170.595 ;
        RECT 311.515 170.510 311.830 171.085 ;
        RECT 311.505 169.845 311.835 170.325 ;
        RECT 312.020 170.125 312.400 171.085 ;
        RECT 312.850 170.755 313.175 171.170 ;
        RECT 313.345 170.755 313.685 171.450 ;
        RECT 313.345 170.585 313.515 170.755 ;
        RECT 313.855 170.585 314.085 172.225 ;
        RECT 314.255 171.425 314.545 172.395 ;
        RECT 314.725 171.305 315.935 172.395 ;
        RECT 312.775 170.415 313.515 170.585 ;
        RECT 312.775 170.015 312.965 170.415 ;
        RECT 313.685 170.395 314.085 170.585 ;
        RECT 314.725 170.595 315.245 171.135 ;
        RECT 315.415 170.765 315.935 171.305 ;
        RECT 316.105 171.305 317.315 172.395 ;
        RECT 316.105 170.765 316.625 171.305 ;
        RECT 316.795 170.595 317.315 171.135 ;
        RECT 313.185 169.845 313.515 170.205 ;
        RECT 313.685 170.015 313.875 170.395 ;
        RECT 314.045 169.845 314.375 170.225 ;
        RECT 314.725 169.845 315.935 170.595 ;
        RECT 316.105 169.845 317.315 170.595 ;
        RECT 388.125 170.375 388.375 173.875 ;
        RECT 389.665 172.750 389.835 173.250 ;
        RECT 388.780 171.480 389.260 172.520 ;
        RECT 389.530 171.480 389.970 172.520 ;
        RECT 390.240 171.480 390.720 172.520 ;
        RECT 389.665 170.750 389.835 171.250 ;
        RECT 391.125 170.375 391.375 173.875 ;
        RECT 388.125 170.125 391.375 170.375 ;
        RECT 293.020 169.675 317.400 169.845 ;
        RECT 293.105 168.925 294.315 169.675 ;
        RECT 294.485 169.130 299.830 169.675 ;
        RECT 300.005 169.130 305.350 169.675 ;
        RECT 305.525 169.130 310.870 169.675 ;
        RECT 293.105 168.385 293.625 168.925 ;
        RECT 293.795 168.215 294.315 168.755 ;
        RECT 296.070 168.300 296.410 169.130 ;
        RECT 293.105 167.125 294.315 168.215 ;
        RECT 297.890 167.560 298.240 168.810 ;
        RECT 301.590 168.300 301.930 169.130 ;
        RECT 303.410 167.560 303.760 168.810 ;
        RECT 307.110 168.300 307.450 169.130 ;
        RECT 311.045 168.925 312.255 169.675 ;
        RECT 312.515 169.125 312.685 169.505 ;
        RECT 312.900 169.295 313.230 169.675 ;
        RECT 312.515 168.955 313.230 169.125 ;
        RECT 308.930 167.560 309.280 168.810 ;
        RECT 311.045 168.385 311.565 168.925 ;
        RECT 311.735 168.215 312.255 168.755 ;
        RECT 312.425 168.405 312.780 168.775 ;
        RECT 313.060 168.765 313.230 168.955 ;
        RECT 313.400 168.930 313.655 169.505 ;
        RECT 313.060 168.435 313.315 168.765 ;
        RECT 313.060 168.225 313.230 168.435 ;
        RECT 294.485 167.125 299.830 167.560 ;
        RECT 300.005 167.125 305.350 167.560 ;
        RECT 305.525 167.125 310.870 167.560 ;
        RECT 311.045 167.125 312.255 168.215 ;
        RECT 312.515 168.055 313.230 168.225 ;
        RECT 313.485 168.200 313.655 168.930 ;
        RECT 313.830 168.835 314.090 169.675 ;
        RECT 314.265 168.905 315.935 169.675 ;
        RECT 316.105 168.925 317.315 169.675 ;
        RECT 314.265 168.385 315.015 168.905 ;
        RECT 312.515 167.295 312.685 168.055 ;
        RECT 312.900 167.125 313.230 167.885 ;
        RECT 313.400 167.295 313.655 168.200 ;
        RECT 313.830 167.125 314.090 168.275 ;
        RECT 315.185 168.215 315.935 168.735 ;
        RECT 314.265 167.125 315.935 168.215 ;
        RECT 316.105 168.215 316.625 168.755 ;
        RECT 316.795 168.385 317.315 168.925 ;
        RECT 316.105 167.125 317.315 168.215 ;
        RECT 293.020 166.955 317.400 167.125 ;
        RECT 293.105 165.865 294.315 166.955 ;
        RECT 294.485 165.865 297.075 166.955 ;
        RECT 297.810 166.495 297.980 166.955 ;
        RECT 298.150 166.325 298.480 166.785 ;
        RECT 293.105 165.155 293.625 165.695 ;
        RECT 293.795 165.325 294.315 165.865 ;
        RECT 294.485 165.175 295.695 165.695 ;
        RECT 295.865 165.345 297.075 165.865 ;
        RECT 297.705 166.155 298.480 166.325 ;
        RECT 298.650 166.155 298.820 166.955 ;
        RECT 293.105 164.405 294.315 165.155 ;
        RECT 294.485 164.405 297.075 165.175 ;
        RECT 297.705 165.145 298.135 166.155 ;
        RECT 299.405 165.985 299.765 166.160 ;
        RECT 298.305 165.815 299.765 165.985 ;
        RECT 300.465 165.945 300.725 166.955 ;
        RECT 300.895 166.115 301.170 166.785 ;
        RECT 298.305 165.315 298.475 165.815 ;
        RECT 297.705 164.975 298.400 165.145 ;
        RECT 298.645 165.085 299.055 165.645 ;
        RECT 297.730 164.405 298.060 164.805 ;
        RECT 298.230 164.705 298.400 164.975 ;
        RECT 299.225 164.915 299.405 165.815 ;
        RECT 300.895 165.765 301.065 166.115 ;
        RECT 301.370 166.110 301.585 166.955 ;
        RECT 301.770 166.445 302.245 166.785 ;
        RECT 302.425 166.450 303.055 166.955 ;
        RECT 302.425 166.275 302.615 166.450 ;
        RECT 301.810 165.915 302.060 166.210 ;
        RECT 302.285 166.085 302.615 166.275 ;
        RECT 302.785 165.915 303.040 166.280 ;
        RECT 299.575 165.255 299.770 165.645 ;
        RECT 299.575 165.085 299.775 165.255 ;
        RECT 300.465 165.245 301.080 165.765 ;
        RECT 301.250 165.745 303.040 165.915 ;
        RECT 303.225 165.865 305.815 166.955 ;
        RECT 301.250 165.315 301.480 165.745 ;
        RECT 298.570 164.405 298.885 164.915 ;
        RECT 299.115 164.575 299.405 164.915 ;
        RECT 299.575 164.405 299.815 164.915 ;
        RECT 300.465 164.405 300.740 165.065 ;
        RECT 300.910 165.035 301.080 165.245 ;
        RECT 301.665 165.070 302.075 165.565 ;
        RECT 300.910 164.575 301.160 165.035 ;
        RECT 301.335 164.405 301.665 164.900 ;
        RECT 301.845 164.625 302.075 165.070 ;
        RECT 302.245 164.890 302.500 165.745 ;
        RECT 302.670 165.085 303.055 165.565 ;
        RECT 303.225 165.175 304.435 165.695 ;
        RECT 304.605 165.345 305.815 165.865 ;
        RECT 305.985 165.790 306.275 166.955 ;
        RECT 306.445 165.865 309.955 166.955 ;
        RECT 310.645 166.255 310.865 166.785 ;
        RECT 311.035 166.445 311.365 166.955 ;
        RECT 311.535 166.255 311.760 166.785 ;
        RECT 310.645 165.990 311.760 166.255 ;
        RECT 311.930 166.240 312.245 166.785 ;
        RECT 312.435 166.540 312.765 166.955 ;
        RECT 311.930 166.010 312.765 166.240 ;
        RECT 306.445 165.175 308.095 165.695 ;
        RECT 308.265 165.345 309.955 165.865 ;
        RECT 302.245 164.625 303.035 164.890 ;
        RECT 303.225 164.405 305.815 165.175 ;
        RECT 305.985 164.405 306.275 165.130 ;
        RECT 306.445 164.405 309.955 165.175 ;
        RECT 310.595 165.070 310.910 165.645 ;
        RECT 310.585 164.405 310.915 164.885 ;
        RECT 311.100 164.685 311.480 165.645 ;
        RECT 311.930 165.315 312.255 165.730 ;
        RECT 312.425 165.315 312.765 166.010 ;
        RECT 312.425 165.145 312.595 165.315 ;
        RECT 312.935 165.145 313.165 166.785 ;
        RECT 313.335 165.985 313.625 166.955 ;
        RECT 313.805 165.865 315.475 166.955 ;
        RECT 311.855 164.975 312.595 165.145 ;
        RECT 311.855 164.575 312.045 164.975 ;
        RECT 312.765 164.955 313.165 165.145 ;
        RECT 313.805 165.175 314.555 165.695 ;
        RECT 314.725 165.345 315.475 165.865 ;
        RECT 316.105 165.865 317.315 166.955 ;
        RECT 388.125 166.625 388.375 170.125 ;
        RECT 389.665 169.000 389.835 169.500 ;
        RECT 388.780 167.730 389.260 168.770 ;
        RECT 389.530 167.730 389.970 168.770 ;
        RECT 390.240 167.730 390.720 168.770 ;
        RECT 389.665 167.000 389.835 167.500 ;
        RECT 391.125 166.625 391.375 170.125 ;
        RECT 388.125 166.375 391.375 166.625 ;
        RECT 397.625 196.375 400.875 196.625 ;
        RECT 397.625 192.875 397.875 196.375 ;
        RECT 399.165 195.250 399.335 195.750 ;
        RECT 398.280 193.980 398.760 195.020 ;
        RECT 399.030 193.980 399.470 195.020 ;
        RECT 399.740 193.980 400.220 195.020 ;
        RECT 399.165 193.250 399.335 193.750 ;
        RECT 400.625 192.875 400.875 196.375 ;
        RECT 397.625 192.625 400.875 192.875 ;
        RECT 397.625 189.125 397.875 192.625 ;
        RECT 399.165 191.500 399.335 192.000 ;
        RECT 398.280 190.230 398.760 191.270 ;
        RECT 399.030 190.230 399.470 191.270 ;
        RECT 399.740 190.230 400.220 191.270 ;
        RECT 399.165 189.500 399.335 190.000 ;
        RECT 400.625 189.125 400.875 192.625 ;
        RECT 397.625 188.875 400.875 189.125 ;
        RECT 397.625 185.375 397.875 188.875 ;
        RECT 399.165 187.750 399.335 188.250 ;
        RECT 398.280 186.480 398.760 187.520 ;
        RECT 399.030 186.480 399.470 187.520 ;
        RECT 399.740 186.480 400.220 187.520 ;
        RECT 399.165 185.750 399.335 186.250 ;
        RECT 400.625 185.375 400.875 188.875 ;
        RECT 397.625 185.125 400.875 185.375 ;
        RECT 397.625 181.625 397.875 185.125 ;
        RECT 399.165 184.000 399.335 184.500 ;
        RECT 398.280 182.730 398.760 183.770 ;
        RECT 399.030 182.730 399.470 183.770 ;
        RECT 399.740 182.730 400.220 183.770 ;
        RECT 399.165 182.000 399.335 182.500 ;
        RECT 400.625 181.625 400.875 185.125 ;
        RECT 397.625 181.375 400.875 181.625 ;
        RECT 397.625 177.875 397.875 181.375 ;
        RECT 399.165 180.250 399.335 180.750 ;
        RECT 398.280 178.980 398.760 180.020 ;
        RECT 399.030 178.980 399.470 180.020 ;
        RECT 399.740 178.980 400.220 180.020 ;
        RECT 399.165 178.250 399.335 178.750 ;
        RECT 400.625 177.875 400.875 181.375 ;
        RECT 397.625 177.625 400.875 177.875 ;
        RECT 397.625 174.125 397.875 177.625 ;
        RECT 399.165 176.500 399.335 177.000 ;
        RECT 398.280 175.230 398.760 176.270 ;
        RECT 399.030 175.230 399.470 176.270 ;
        RECT 399.740 175.230 400.220 176.270 ;
        RECT 399.165 174.500 399.335 175.000 ;
        RECT 400.625 174.125 400.875 177.625 ;
        RECT 397.625 173.875 400.875 174.125 ;
        RECT 397.625 170.375 397.875 173.875 ;
        RECT 399.165 172.750 399.335 173.250 ;
        RECT 398.280 171.480 398.760 172.520 ;
        RECT 399.030 171.480 399.470 172.520 ;
        RECT 399.740 171.480 400.220 172.520 ;
        RECT 399.165 170.750 399.335 171.250 ;
        RECT 400.625 170.375 400.875 173.875 ;
        RECT 397.625 170.125 400.875 170.375 ;
        RECT 397.625 166.625 397.875 170.125 ;
        RECT 399.165 169.000 399.335 169.500 ;
        RECT 398.280 167.730 398.760 168.770 ;
        RECT 399.030 167.730 399.470 168.770 ;
        RECT 399.740 167.730 400.220 168.770 ;
        RECT 399.165 167.000 399.335 167.500 ;
        RECT 400.625 166.625 400.875 170.125 ;
        RECT 397.625 166.375 400.875 166.625 ;
        RECT 407.125 196.375 410.375 196.625 ;
        RECT 407.125 192.875 407.375 196.375 ;
        RECT 408.665 195.250 408.835 195.750 ;
        RECT 407.780 193.980 408.260 195.020 ;
        RECT 408.530 193.980 408.970 195.020 ;
        RECT 409.240 193.980 409.720 195.020 ;
        RECT 408.665 193.250 408.835 193.750 ;
        RECT 410.125 192.875 410.375 196.375 ;
        RECT 407.125 192.625 410.375 192.875 ;
        RECT 407.125 189.125 407.375 192.625 ;
        RECT 408.665 191.500 408.835 192.000 ;
        RECT 407.780 190.230 408.260 191.270 ;
        RECT 408.530 190.230 408.970 191.270 ;
        RECT 409.240 190.230 409.720 191.270 ;
        RECT 408.665 189.500 408.835 190.000 ;
        RECT 410.125 189.125 410.375 192.625 ;
        RECT 407.125 188.875 410.375 189.125 ;
        RECT 407.125 185.375 407.375 188.875 ;
        RECT 408.665 187.750 408.835 188.250 ;
        RECT 407.780 186.480 408.260 187.520 ;
        RECT 408.530 186.480 408.970 187.520 ;
        RECT 409.240 186.480 409.720 187.520 ;
        RECT 408.665 185.750 408.835 186.250 ;
        RECT 410.125 185.375 410.375 188.875 ;
        RECT 407.125 185.125 410.375 185.375 ;
        RECT 407.125 181.625 407.375 185.125 ;
        RECT 408.665 184.000 408.835 184.500 ;
        RECT 407.780 182.730 408.260 183.770 ;
        RECT 408.530 182.730 408.970 183.770 ;
        RECT 409.240 182.730 409.720 183.770 ;
        RECT 408.665 182.000 408.835 182.500 ;
        RECT 410.125 181.625 410.375 185.125 ;
        RECT 407.125 181.375 410.375 181.625 ;
        RECT 407.125 177.875 407.375 181.375 ;
        RECT 408.665 180.250 408.835 180.750 ;
        RECT 407.780 178.980 408.260 180.020 ;
        RECT 408.530 178.980 408.970 180.020 ;
        RECT 409.240 178.980 409.720 180.020 ;
        RECT 408.665 178.250 408.835 178.750 ;
        RECT 410.125 177.875 410.375 181.375 ;
        RECT 407.125 177.625 410.375 177.875 ;
        RECT 407.125 174.125 407.375 177.625 ;
        RECT 408.665 176.500 408.835 177.000 ;
        RECT 407.780 175.230 408.260 176.270 ;
        RECT 408.530 175.230 408.970 176.270 ;
        RECT 409.240 175.230 409.720 176.270 ;
        RECT 408.665 174.500 408.835 175.000 ;
        RECT 410.125 174.125 410.375 177.625 ;
        RECT 407.125 173.875 410.375 174.125 ;
        RECT 407.125 170.375 407.375 173.875 ;
        RECT 408.665 172.750 408.835 173.250 ;
        RECT 407.780 171.480 408.260 172.520 ;
        RECT 408.530 171.480 408.970 172.520 ;
        RECT 409.240 171.480 409.720 172.520 ;
        RECT 408.665 170.750 408.835 171.250 ;
        RECT 410.125 170.375 410.375 173.875 ;
        RECT 407.125 170.125 410.375 170.375 ;
        RECT 407.125 166.625 407.375 170.125 ;
        RECT 408.665 169.000 408.835 169.500 ;
        RECT 407.780 167.730 408.260 168.770 ;
        RECT 408.530 167.730 408.970 168.770 ;
        RECT 409.240 167.730 409.720 168.770 ;
        RECT 408.665 167.000 408.835 167.500 ;
        RECT 410.125 166.625 410.375 170.125 ;
        RECT 407.125 166.375 410.375 166.625 ;
        RECT 316.105 165.325 316.625 165.865 ;
        RECT 312.265 164.405 312.595 164.765 ;
        RECT 312.765 164.575 312.955 164.955 ;
        RECT 313.125 164.405 313.455 164.785 ;
        RECT 313.805 164.405 315.475 165.175 ;
        RECT 316.795 165.155 317.315 165.695 ;
        RECT 316.105 164.405 317.315 165.155 ;
        RECT 390.875 165.125 409.125 165.375 ;
        RECT 293.020 164.235 317.400 164.405 ;
        RECT 293.105 163.485 294.315 164.235 ;
        RECT 294.665 163.575 295.005 164.235 ;
        RECT 293.105 162.945 293.625 163.485 ;
        RECT 293.795 162.775 294.315 163.315 ;
        RECT 293.105 161.685 294.315 162.775 ;
        RECT 294.485 161.855 295.005 163.405 ;
        RECT 295.175 162.580 295.695 164.065 ;
        RECT 296.045 163.855 296.375 164.235 ;
        RECT 296.545 163.685 296.735 164.065 ;
        RECT 296.905 163.875 297.235 164.235 ;
        RECT 296.335 163.495 296.735 163.685 ;
        RECT 297.455 163.665 297.645 164.065 ;
        RECT 296.905 163.495 297.645 163.665 ;
        RECT 295.175 161.685 295.505 162.410 ;
        RECT 295.875 161.685 296.165 162.655 ;
        RECT 296.335 161.855 296.565 163.495 ;
        RECT 296.905 163.325 297.075 163.495 ;
        RECT 296.735 162.630 297.075 163.325 ;
        RECT 297.245 162.910 297.570 163.325 ;
        RECT 298.020 162.995 298.400 163.955 ;
        RECT 298.585 163.755 298.915 164.235 ;
        RECT 298.590 162.995 298.905 163.570 ;
        RECT 299.085 163.435 299.375 164.235 ;
        RECT 299.545 163.775 300.095 164.065 ;
        RECT 300.265 163.775 300.515 164.235 ;
        RECT 296.735 162.400 297.570 162.630 ;
        RECT 296.735 161.685 297.065 162.100 ;
        RECT 297.255 161.855 297.570 162.400 ;
        RECT 297.740 162.385 298.855 162.650 ;
        RECT 297.740 161.855 297.965 162.385 ;
        RECT 298.135 161.685 298.465 162.195 ;
        RECT 298.635 161.855 298.855 162.385 ;
        RECT 299.085 161.685 299.375 162.825 ;
        RECT 299.545 162.405 299.795 163.775 ;
        RECT 301.145 163.605 301.475 163.965 ;
        RECT 301.845 163.690 307.190 164.235 ;
        RECT 300.085 163.415 301.475 163.605 ;
        RECT 300.085 163.325 300.255 163.415 ;
        RECT 299.965 162.995 300.255 163.325 ;
        RECT 300.425 162.995 300.755 163.245 ;
        RECT 300.985 162.995 301.675 163.245 ;
        RECT 300.085 162.745 300.255 162.995 ;
        RECT 300.085 162.575 301.025 162.745 ;
        RECT 299.545 161.855 299.995 162.405 ;
        RECT 300.185 161.685 300.515 162.405 ;
        RECT 300.725 162.025 301.025 162.575 ;
        RECT 301.360 162.555 301.675 162.995 ;
        RECT 303.430 162.860 303.770 163.690 ;
        RECT 307.365 163.465 310.875 164.235 ;
        RECT 311.505 163.755 311.835 164.235 ;
        RECT 301.195 161.685 301.475 162.355 ;
        RECT 305.250 162.120 305.600 163.370 ;
        RECT 307.365 162.945 309.015 163.465 ;
        RECT 309.185 162.775 310.875 163.295 ;
        RECT 311.515 162.995 311.830 163.570 ;
        RECT 312.020 162.995 312.400 163.955 ;
        RECT 312.775 163.665 312.965 164.065 ;
        RECT 313.185 163.875 313.515 164.235 ;
        RECT 313.685 163.685 313.875 164.065 ;
        RECT 314.045 163.855 314.375 164.235 ;
        RECT 312.775 163.495 313.515 163.665 ;
        RECT 313.685 163.495 314.085 163.685 ;
        RECT 313.345 163.325 313.515 163.495 ;
        RECT 312.850 162.910 313.175 163.325 ;
        RECT 301.845 161.685 307.190 162.120 ;
        RECT 307.365 161.685 310.875 162.775 ;
        RECT 311.565 162.385 312.680 162.650 ;
        RECT 313.345 162.630 313.685 163.325 ;
        RECT 311.565 161.855 311.785 162.385 ;
        RECT 311.955 161.685 312.285 162.195 ;
        RECT 312.455 161.855 312.680 162.385 ;
        RECT 312.850 162.400 313.685 162.630 ;
        RECT 312.850 161.855 313.165 162.400 ;
        RECT 313.355 161.685 313.685 162.100 ;
        RECT 313.855 161.855 314.085 163.495 ;
        RECT 314.725 163.485 315.935 164.235 ;
        RECT 316.105 163.485 317.315 164.235 ;
        RECT 314.725 162.945 315.245 163.485 ;
        RECT 315.415 162.775 315.935 163.315 ;
        RECT 314.255 161.685 314.545 162.655 ;
        RECT 314.725 161.685 315.935 162.775 ;
        RECT 316.105 162.775 316.625 163.315 ;
        RECT 316.795 162.945 317.315 163.485 ;
        RECT 379.375 163.625 390.125 163.875 ;
        RECT 316.105 161.685 317.315 162.775 ;
        RECT 293.020 161.515 317.400 161.685 ;
        RECT 293.105 160.425 294.315 161.515 ;
        RECT 294.485 161.080 299.830 161.515 ;
        RECT 300.005 161.080 305.350 161.515 ;
        RECT 293.105 159.715 293.625 160.255 ;
        RECT 293.795 159.885 294.315 160.425 ;
        RECT 293.105 158.965 294.315 159.715 ;
        RECT 296.070 159.510 296.410 160.340 ;
        RECT 297.890 159.830 298.240 161.080 ;
        RECT 301.590 159.510 301.930 160.340 ;
        RECT 303.410 159.830 303.760 161.080 ;
        RECT 305.985 160.350 306.275 161.515 ;
        RECT 306.445 161.080 311.790 161.515 ;
        RECT 294.485 158.965 299.830 159.510 ;
        RECT 300.005 158.965 305.350 159.510 ;
        RECT 305.985 158.965 306.275 159.690 ;
        RECT 308.030 159.510 308.370 160.340 ;
        RECT 309.850 159.830 310.200 161.080 ;
        RECT 311.965 160.425 315.475 161.515 ;
        RECT 311.965 159.735 313.615 160.255 ;
        RECT 313.785 159.905 315.475 160.425 ;
        RECT 316.105 160.425 317.315 161.515 ;
        RECT 316.105 159.885 316.625 160.425 ;
        RECT 306.445 158.965 311.790 159.510 ;
        RECT 311.965 158.965 315.475 159.735 ;
        RECT 316.795 159.715 317.315 160.255 ;
        RECT 316.105 158.965 317.315 159.715 ;
        RECT 293.020 158.795 317.400 158.965 ;
        RECT 379.375 152.875 379.625 163.625 ;
        RECT 380.915 162.750 381.585 163.250 ;
        RECT 380.030 153.980 380.690 162.520 ;
        RECT 381.810 153.980 382.470 162.520 ;
        RECT 380.915 153.250 381.585 153.750 ;
        RECT 382.875 152.875 383.125 163.625 ;
        RECT 384.415 162.750 385.085 163.250 ;
        RECT 383.530 153.980 384.190 162.520 ;
        RECT 385.310 153.980 385.970 162.520 ;
        RECT 384.415 153.250 385.085 153.750 ;
        RECT 386.375 152.875 386.625 163.625 ;
        RECT 387.915 162.750 388.585 163.250 ;
        RECT 387.030 153.980 387.690 162.520 ;
        RECT 388.810 153.980 389.470 162.520 ;
        RECT 387.915 153.250 388.585 153.750 ;
        RECT 389.875 152.875 390.125 163.625 ;
        RECT 390.875 158.875 391.125 165.125 ;
        RECT 391.615 160.730 391.785 164.770 ;
        RECT 392.075 160.730 392.245 164.770 ;
        RECT 392.535 160.730 392.705 164.770 ;
        RECT 392.995 160.730 393.165 164.770 ;
        RECT 393.455 160.730 393.625 164.770 ;
        RECT 393.915 160.730 394.085 164.770 ;
        RECT 394.375 160.730 394.545 164.770 ;
        RECT 394.835 160.730 395.005 164.770 ;
        RECT 395.295 160.730 395.465 164.770 ;
        RECT 395.755 160.730 395.925 164.770 ;
        RECT 396.215 160.730 396.385 164.770 ;
        RECT 393.915 159.250 394.085 159.750 ;
        RECT 396.875 158.875 397.125 165.125 ;
        RECT 397.615 160.730 397.785 164.770 ;
        RECT 398.075 160.730 398.245 164.770 ;
        RECT 398.535 160.730 398.705 164.770 ;
        RECT 398.995 160.730 399.165 164.770 ;
        RECT 399.455 160.730 399.625 164.770 ;
        RECT 399.915 160.730 400.085 164.770 ;
        RECT 400.375 160.730 400.545 164.770 ;
        RECT 400.835 160.730 401.005 164.770 ;
        RECT 401.295 160.730 401.465 164.770 ;
        RECT 401.755 160.730 401.925 164.770 ;
        RECT 402.215 160.730 402.385 164.770 ;
        RECT 399.915 159.250 400.085 159.750 ;
        RECT 402.875 158.875 403.125 165.125 ;
        RECT 403.615 160.730 403.785 164.770 ;
        RECT 404.075 160.730 404.245 164.770 ;
        RECT 404.535 160.730 404.705 164.770 ;
        RECT 404.995 160.730 405.165 164.770 ;
        RECT 405.455 160.730 405.625 164.770 ;
        RECT 405.915 160.730 406.085 164.770 ;
        RECT 406.375 160.730 406.545 164.770 ;
        RECT 406.835 160.730 407.005 164.770 ;
        RECT 407.295 160.730 407.465 164.770 ;
        RECT 407.755 160.730 407.925 164.770 ;
        RECT 408.215 160.730 408.385 164.770 ;
        RECT 405.915 159.250 406.085 159.750 ;
        RECT 408.875 158.875 409.125 165.125 ;
        RECT 390.875 158.625 409.125 158.875 ;
        RECT 409.625 163.125 420.875 163.375 ;
        RECT 409.625 158.875 409.875 163.125 ;
        RECT 410.215 160.730 410.385 162.770 ;
        RECT 410.655 160.730 410.825 162.770 ;
        RECT 411.095 160.730 411.265 162.770 ;
        RECT 411.535 160.730 411.705 162.770 ;
        RECT 411.975 160.730 412.145 162.770 ;
        RECT 412.415 160.730 412.585 162.770 ;
        RECT 412.855 160.730 413.025 162.770 ;
        RECT 413.295 160.730 413.465 162.770 ;
        RECT 413.735 160.730 413.905 162.770 ;
        RECT 414.175 160.730 414.345 162.770 ;
        RECT 414.615 160.730 414.785 162.770 ;
        RECT 412.420 159.250 412.590 159.750 ;
        RECT 415.125 158.875 415.375 163.125 ;
        RECT 415.715 160.730 415.885 162.770 ;
        RECT 416.155 160.730 416.325 162.770 ;
        RECT 416.595 160.730 416.765 162.770 ;
        RECT 417.035 160.730 417.205 162.770 ;
        RECT 417.475 160.730 417.645 162.770 ;
        RECT 417.915 160.730 418.085 162.770 ;
        RECT 418.355 160.730 418.525 162.770 ;
        RECT 418.795 160.730 418.965 162.770 ;
        RECT 419.235 160.730 419.405 162.770 ;
        RECT 419.675 160.730 419.845 162.770 ;
        RECT 420.115 160.730 420.285 162.770 ;
        RECT 417.920 159.250 418.090 159.750 ;
        RECT 420.625 158.875 420.875 163.125 ;
        RECT 409.625 158.625 420.875 158.875 ;
        RECT 379.375 152.625 390.125 152.875 ;
        RECT 390.875 157.625 409.125 157.875 ;
        RECT 286.250 151.250 354.500 151.750 ;
        RECT 286.250 127.250 286.750 151.250 ;
        RECT 287.250 148.125 344.500 148.375 ;
        RECT 287.430 146.535 287.820 148.125 ;
        RECT 288.030 147.000 288.200 147.830 ;
        RECT 288.570 147.630 288.900 147.800 ;
        RECT 288.030 146.500 288.320 147.000 ;
        RECT 287.430 144.365 287.820 145.730 ;
        RECT 288.030 144.685 288.200 146.500 ;
        RECT 288.490 146.475 288.880 147.415 ;
        RECT 289.330 146.475 289.500 148.125 ;
        RECT 289.830 147.630 290.160 147.800 ;
        RECT 289.890 146.475 290.160 147.415 ;
        RECT 290.330 146.475 290.500 148.125 ;
        RECT 288.370 145.855 288.540 146.185 ;
        RECT 288.710 146.105 288.880 146.475 ;
        RECT 289.990 146.185 290.160 146.475 ;
        RECT 290.770 146.185 290.940 147.415 ;
        RECT 291.330 146.475 291.500 148.125 ;
        RECT 291.770 146.475 292.040 147.415 ;
        RECT 292.210 146.475 292.380 148.125 ;
        RECT 293.030 147.000 293.200 147.830 ;
        RECT 293.570 147.630 293.900 147.800 ;
        RECT 293.030 146.500 293.320 147.000 ;
        RECT 288.710 145.935 289.820 146.105 ;
        RECT 288.710 145.565 288.880 145.935 ;
        RECT 289.990 145.860 290.600 146.185 ;
        RECT 289.990 145.565 290.160 145.860 ;
        RECT 290.430 145.855 290.600 145.860 ;
        RECT 290.770 145.855 291.700 146.185 ;
        RECT 290.770 145.565 290.940 145.855 ;
        RECT 291.870 145.565 292.040 146.475 ;
        RECT 288.610 145.075 288.880 145.565 ;
        RECT 289.050 144.365 289.220 145.565 ;
        RECT 289.890 145.075 290.160 145.565 ;
        RECT 290.490 145.395 290.940 145.565 ;
        RECT 290.490 145.075 290.660 145.395 ;
        RECT 289.390 144.535 290.900 144.885 ;
        RECT 291.330 144.365 291.500 145.565 ;
        RECT 291.770 145.075 292.040 145.565 ;
        RECT 292.210 144.365 292.380 145.565 ;
        RECT 293.030 144.685 293.200 146.500 ;
        RECT 293.490 146.475 293.880 147.415 ;
        RECT 294.330 146.475 294.500 148.125 ;
        RECT 294.830 147.630 295.160 147.800 ;
        RECT 294.890 146.475 295.160 147.415 ;
        RECT 295.330 146.475 295.500 148.125 ;
        RECT 293.370 145.855 293.540 146.185 ;
        RECT 293.710 146.105 293.880 146.475 ;
        RECT 294.990 146.185 295.160 146.475 ;
        RECT 295.770 146.185 295.940 147.415 ;
        RECT 296.330 146.475 296.500 148.125 ;
        RECT 296.770 146.475 297.040 147.415 ;
        RECT 297.210 146.475 297.380 148.125 ;
        RECT 298.115 146.475 298.285 148.125 ;
        RECT 298.555 146.475 298.725 147.415 ;
        RECT 298.995 146.475 299.165 148.125 ;
        RECT 299.850 146.475 300.020 148.125 ;
        RECT 300.690 146.475 300.860 147.415 ;
        RECT 301.430 146.535 301.820 148.125 ;
        RECT 302.350 146.475 302.520 148.125 ;
        RECT 303.190 146.475 303.360 147.415 ;
        RECT 304.030 147.000 304.200 147.830 ;
        RECT 304.570 147.630 304.900 147.800 ;
        RECT 304.030 146.500 304.320 147.000 ;
        RECT 293.710 145.935 294.820 146.105 ;
        RECT 293.710 145.565 293.880 145.935 ;
        RECT 294.990 145.860 295.600 146.185 ;
        RECT 294.990 145.565 295.160 145.860 ;
        RECT 295.430 145.855 295.600 145.860 ;
        RECT 295.770 145.855 296.700 146.185 ;
        RECT 295.770 145.565 295.940 145.855 ;
        RECT 296.870 145.565 297.040 146.475 ;
        RECT 298.030 146.185 298.885 146.265 ;
        RECT 298.000 145.855 298.885 146.185 ;
        RECT 299.750 146.090 300.080 146.305 ;
        RECT 300.250 146.135 300.940 146.305 ;
        RECT 298.030 145.775 298.885 145.855 ;
        RECT 293.610 145.075 293.880 145.565 ;
        RECT 294.050 144.365 294.220 145.565 ;
        RECT 294.890 145.075 295.160 145.565 ;
        RECT 295.490 145.395 295.940 145.565 ;
        RECT 295.490 145.075 295.660 145.395 ;
        RECT 294.390 144.535 295.900 144.885 ;
        RECT 296.330 144.365 296.500 145.565 ;
        RECT 296.770 145.075 297.040 145.565 ;
        RECT 297.210 144.365 297.380 145.565 ;
        RECT 298.115 144.365 298.285 145.565 ;
        RECT 298.555 145.075 298.725 145.565 ;
        RECT 298.995 144.365 299.165 145.565 ;
        RECT 299.810 144.365 299.980 145.565 ;
        RECT 300.250 145.075 300.420 146.135 ;
        RECT 302.250 146.090 302.580 146.305 ;
        RECT 302.750 146.135 303.440 146.305 ;
        RECT 300.590 145.735 300.920 145.905 ;
        RECT 300.690 144.365 300.860 145.565 ;
        RECT 301.430 144.365 301.820 145.730 ;
        RECT 302.310 144.365 302.480 145.565 ;
        RECT 302.750 145.075 302.920 146.135 ;
        RECT 303.090 145.735 303.420 145.905 ;
        RECT 303.190 144.365 303.360 145.565 ;
        RECT 304.030 144.685 304.200 146.500 ;
        RECT 304.490 146.475 304.880 147.415 ;
        RECT 305.330 146.475 305.500 148.125 ;
        RECT 305.830 147.630 306.160 147.800 ;
        RECT 305.890 146.475 306.160 147.415 ;
        RECT 306.330 146.475 306.500 148.125 ;
        RECT 304.370 145.855 304.540 146.185 ;
        RECT 304.710 146.105 304.880 146.475 ;
        RECT 305.990 146.185 306.160 146.475 ;
        RECT 306.770 146.185 306.940 147.415 ;
        RECT 307.330 146.475 307.500 148.125 ;
        RECT 307.770 146.475 308.040 147.415 ;
        RECT 308.210 146.475 308.380 148.125 ;
        RECT 309.030 147.000 309.200 147.830 ;
        RECT 309.570 147.630 309.900 147.800 ;
        RECT 309.030 146.500 309.320 147.000 ;
        RECT 304.710 145.935 305.820 146.105 ;
        RECT 304.710 145.565 304.880 145.935 ;
        RECT 305.990 145.860 306.600 146.185 ;
        RECT 305.990 145.565 306.160 145.860 ;
        RECT 306.430 145.855 306.600 145.860 ;
        RECT 306.770 145.855 307.700 146.185 ;
        RECT 306.770 145.565 306.940 145.855 ;
        RECT 307.870 145.565 308.040 146.475 ;
        RECT 304.610 145.075 304.880 145.565 ;
        RECT 305.050 144.365 305.220 145.565 ;
        RECT 305.890 145.075 306.160 145.565 ;
        RECT 306.490 145.395 306.940 145.565 ;
        RECT 306.490 145.075 306.660 145.395 ;
        RECT 305.390 144.535 306.900 144.885 ;
        RECT 307.330 144.365 307.500 145.565 ;
        RECT 307.770 145.075 308.040 145.565 ;
        RECT 308.210 144.365 308.380 145.565 ;
        RECT 309.030 144.685 309.200 146.500 ;
        RECT 309.490 146.475 309.880 147.415 ;
        RECT 310.330 146.475 310.500 148.125 ;
        RECT 310.830 147.630 311.160 147.800 ;
        RECT 310.890 146.475 311.160 147.415 ;
        RECT 311.330 146.475 311.500 148.125 ;
        RECT 309.370 145.855 309.540 146.185 ;
        RECT 309.710 146.105 309.880 146.475 ;
        RECT 310.990 146.185 311.160 146.475 ;
        RECT 311.770 146.185 311.940 147.415 ;
        RECT 312.330 146.475 312.500 148.125 ;
        RECT 312.770 146.475 313.040 147.415 ;
        RECT 313.210 146.475 313.380 148.125 ;
        RECT 313.930 146.535 314.320 148.125 ;
        RECT 314.880 146.475 315.050 148.125 ;
        RECT 315.320 146.475 315.590 147.415 ;
        RECT 315.760 146.475 315.930 148.125 ;
        RECT 316.200 146.475 316.370 147.415 ;
        RECT 316.640 146.475 316.810 148.125 ;
        RECT 317.280 147.000 317.450 147.830 ;
        RECT 317.820 147.630 318.150 147.800 ;
        RECT 317.280 146.500 317.570 147.000 ;
        RECT 309.710 145.935 310.820 146.105 ;
        RECT 309.710 145.565 309.880 145.935 ;
        RECT 310.990 145.860 311.600 146.185 ;
        RECT 310.990 145.565 311.160 145.860 ;
        RECT 311.430 145.855 311.600 145.860 ;
        RECT 311.770 145.855 312.700 146.185 ;
        RECT 311.770 145.565 311.940 145.855 ;
        RECT 312.870 145.565 313.040 146.475 ;
        RECT 314.750 146.090 315.290 146.305 ;
        RECT 315.630 146.095 316.320 146.265 ;
        RECT 315.990 146.050 316.320 146.095 ;
        RECT 315.480 145.905 315.810 145.925 ;
        RECT 314.810 145.735 315.810 145.905 ;
        RECT 309.610 145.075 309.880 145.565 ;
        RECT 310.050 144.365 310.220 145.565 ;
        RECT 310.890 145.075 311.160 145.565 ;
        RECT 311.490 145.395 311.940 145.565 ;
        RECT 311.490 145.075 311.660 145.395 ;
        RECT 310.390 144.535 311.900 144.885 ;
        RECT 312.330 144.365 312.500 145.565 ;
        RECT 312.770 145.075 313.040 145.565 ;
        RECT 313.210 144.365 313.380 145.565 ;
        RECT 313.930 144.365 314.320 145.730 ;
        RECT 314.920 145.075 315.590 145.565 ;
        RECT 315.760 144.365 315.930 145.565 ;
        RECT 316.200 145.075 316.370 145.565 ;
        RECT 316.640 144.365 316.810 145.565 ;
        RECT 317.280 144.685 317.450 146.500 ;
        RECT 317.740 146.475 318.130 147.415 ;
        RECT 318.580 146.475 318.750 148.125 ;
        RECT 319.080 147.630 319.410 147.800 ;
        RECT 319.140 146.475 319.410 147.415 ;
        RECT 319.580 146.475 319.750 148.125 ;
        RECT 317.620 145.855 317.790 146.185 ;
        RECT 317.960 146.105 318.130 146.475 ;
        RECT 319.240 146.185 319.410 146.475 ;
        RECT 320.020 146.185 320.190 147.415 ;
        RECT 320.580 146.475 320.750 148.125 ;
        RECT 321.020 146.475 321.290 147.415 ;
        RECT 321.460 146.475 321.630 148.125 ;
        RECT 322.365 146.475 322.535 148.125 ;
        RECT 322.805 146.475 322.975 147.415 ;
        RECT 323.245 146.475 323.415 148.125 ;
        RECT 323.930 146.535 324.320 148.125 ;
        RECT 324.780 147.000 324.950 147.830 ;
        RECT 325.320 147.630 325.650 147.800 ;
        RECT 324.780 146.500 325.070 147.000 ;
        RECT 317.960 145.935 319.070 146.105 ;
        RECT 317.960 145.565 318.130 145.935 ;
        RECT 319.240 145.860 319.850 146.185 ;
        RECT 319.240 145.565 319.410 145.860 ;
        RECT 319.680 145.855 319.850 145.860 ;
        RECT 320.020 145.855 320.950 146.185 ;
        RECT 320.020 145.565 320.190 145.855 ;
        RECT 321.120 145.565 321.290 146.475 ;
        RECT 322.280 146.185 323.135 146.265 ;
        RECT 322.250 145.855 323.135 146.185 ;
        RECT 322.280 145.775 323.135 145.855 ;
        RECT 317.860 145.075 318.130 145.565 ;
        RECT 318.300 144.365 318.470 145.565 ;
        RECT 319.140 145.075 319.410 145.565 ;
        RECT 319.740 145.395 320.190 145.565 ;
        RECT 319.740 145.075 319.910 145.395 ;
        RECT 318.640 144.535 320.150 144.885 ;
        RECT 320.580 144.365 320.750 145.565 ;
        RECT 321.020 145.075 321.290 145.565 ;
        RECT 321.460 144.365 321.630 145.565 ;
        RECT 322.365 144.365 322.535 145.565 ;
        RECT 322.805 145.075 322.975 145.565 ;
        RECT 323.245 144.365 323.415 145.565 ;
        RECT 323.930 144.365 324.320 145.730 ;
        RECT 324.780 144.685 324.950 146.500 ;
        RECT 325.240 146.475 325.630 147.415 ;
        RECT 326.080 146.475 326.250 148.125 ;
        RECT 326.580 147.630 326.910 147.800 ;
        RECT 326.640 146.475 326.910 147.415 ;
        RECT 327.080 146.475 327.250 148.125 ;
        RECT 325.120 145.855 325.290 146.185 ;
        RECT 325.460 146.105 325.630 146.475 ;
        RECT 326.740 146.185 326.910 146.475 ;
        RECT 327.520 146.185 327.690 147.415 ;
        RECT 328.080 146.475 328.250 148.125 ;
        RECT 328.520 146.475 328.790 147.415 ;
        RECT 328.960 146.475 329.130 148.125 ;
        RECT 329.780 147.000 329.950 147.830 ;
        RECT 330.320 147.630 330.650 147.800 ;
        RECT 329.780 146.500 330.070 147.000 ;
        RECT 325.460 145.935 326.570 146.105 ;
        RECT 325.460 145.565 325.630 145.935 ;
        RECT 326.740 145.860 327.350 146.185 ;
        RECT 326.740 145.565 326.910 145.860 ;
        RECT 327.180 145.855 327.350 145.860 ;
        RECT 327.520 145.855 328.450 146.185 ;
        RECT 327.520 145.565 327.690 145.855 ;
        RECT 328.620 145.565 328.790 146.475 ;
        RECT 325.360 145.075 325.630 145.565 ;
        RECT 325.800 144.365 325.970 145.565 ;
        RECT 326.640 145.075 326.910 145.565 ;
        RECT 327.240 145.395 327.690 145.565 ;
        RECT 327.240 145.075 327.410 145.395 ;
        RECT 326.140 144.535 327.650 144.885 ;
        RECT 328.080 144.365 328.250 145.565 ;
        RECT 328.520 145.075 328.790 145.565 ;
        RECT 328.960 144.365 329.130 145.565 ;
        RECT 329.780 144.685 329.950 146.500 ;
        RECT 330.240 146.475 330.630 147.415 ;
        RECT 331.080 146.475 331.250 148.125 ;
        RECT 331.580 147.630 331.910 147.800 ;
        RECT 331.640 146.475 331.910 147.415 ;
        RECT 332.080 146.475 332.250 148.125 ;
        RECT 330.120 145.855 330.290 146.185 ;
        RECT 330.460 146.105 330.630 146.475 ;
        RECT 331.740 146.185 331.910 146.475 ;
        RECT 332.520 146.185 332.690 147.415 ;
        RECT 333.080 146.475 333.250 148.125 ;
        RECT 333.520 146.475 333.790 147.415 ;
        RECT 333.960 146.475 334.130 148.125 ;
        RECT 334.680 146.535 335.070 148.125 ;
        RECT 335.530 147.000 335.700 147.830 ;
        RECT 336.070 147.630 336.400 147.800 ;
        RECT 335.530 146.500 335.820 147.000 ;
        RECT 330.460 145.935 331.570 146.105 ;
        RECT 330.460 145.565 330.630 145.935 ;
        RECT 331.740 145.860 332.350 146.185 ;
        RECT 331.740 145.565 331.910 145.860 ;
        RECT 332.180 145.855 332.350 145.860 ;
        RECT 332.520 145.855 333.450 146.185 ;
        RECT 332.520 145.565 332.690 145.855 ;
        RECT 333.620 145.565 333.790 146.475 ;
        RECT 330.360 145.075 330.630 145.565 ;
        RECT 330.800 144.365 330.970 145.565 ;
        RECT 331.640 145.075 331.910 145.565 ;
        RECT 332.240 145.395 332.690 145.565 ;
        RECT 332.240 145.075 332.410 145.395 ;
        RECT 331.140 144.535 332.650 144.885 ;
        RECT 333.080 144.365 333.250 145.565 ;
        RECT 333.520 145.075 333.790 145.565 ;
        RECT 333.960 144.365 334.130 145.565 ;
        RECT 334.680 144.365 335.070 145.730 ;
        RECT 335.530 144.685 335.700 146.500 ;
        RECT 335.990 146.475 336.380 147.415 ;
        RECT 336.830 146.475 337.000 148.125 ;
        RECT 337.330 147.630 337.660 147.800 ;
        RECT 337.390 146.475 337.660 147.415 ;
        RECT 337.830 146.475 338.000 148.125 ;
        RECT 335.870 145.855 336.040 146.185 ;
        RECT 336.210 146.105 336.380 146.475 ;
        RECT 337.490 146.185 337.660 146.475 ;
        RECT 338.270 146.185 338.440 147.415 ;
        RECT 338.830 146.475 339.000 148.125 ;
        RECT 339.270 146.475 339.540 147.415 ;
        RECT 339.710 146.475 339.880 148.125 ;
        RECT 340.615 146.475 340.785 148.125 ;
        RECT 341.055 146.475 341.225 147.415 ;
        RECT 341.495 146.475 341.665 148.125 ;
        RECT 342.365 146.475 342.535 148.125 ;
        RECT 342.805 146.475 342.975 147.415 ;
        RECT 343.245 146.475 343.415 148.125 ;
        RECT 343.930 146.535 344.320 148.125 ;
        RECT 336.210 145.935 337.320 146.105 ;
        RECT 336.210 145.565 336.380 145.935 ;
        RECT 337.490 145.860 338.100 146.185 ;
        RECT 337.490 145.565 337.660 145.860 ;
        RECT 337.930 145.855 338.100 145.860 ;
        RECT 338.270 145.855 339.200 146.185 ;
        RECT 338.270 145.565 338.440 145.855 ;
        RECT 339.370 145.565 339.540 146.475 ;
        RECT 340.530 146.185 341.385 146.265 ;
        RECT 342.280 146.185 343.135 146.265 ;
        RECT 340.500 145.855 341.385 146.185 ;
        RECT 342.250 145.855 343.135 146.185 ;
        RECT 340.530 145.775 341.385 145.855 ;
        RECT 342.280 145.775 343.135 145.855 ;
        RECT 336.110 145.075 336.380 145.565 ;
        RECT 336.550 144.365 336.720 145.565 ;
        RECT 337.390 145.075 337.660 145.565 ;
        RECT 337.990 145.395 338.440 145.565 ;
        RECT 337.990 145.075 338.160 145.395 ;
        RECT 336.890 144.535 338.400 144.885 ;
        RECT 338.830 144.365 339.000 145.565 ;
        RECT 339.270 145.075 339.540 145.565 ;
        RECT 339.710 144.365 339.880 145.565 ;
        RECT 340.615 144.365 340.785 145.565 ;
        RECT 341.055 145.075 341.225 145.565 ;
        RECT 341.495 144.365 341.665 145.565 ;
        RECT 342.365 144.365 342.535 145.565 ;
        RECT 342.805 145.075 342.975 145.565 ;
        RECT 343.245 144.365 343.415 145.565 ;
        RECT 343.930 144.365 344.320 145.730 ;
        RECT 287.250 144.115 344.500 144.365 ;
        RECT 293.000 141.125 341.250 141.375 ;
        RECT 343.500 141.125 351.000 141.375 ;
        RECT 293.180 139.535 293.570 141.125 ;
        RECT 294.085 139.475 294.255 141.125 ;
        RECT 294.525 139.475 294.695 140.415 ;
        RECT 294.965 139.475 295.135 141.125 ;
        RECT 295.760 139.475 295.930 141.125 ;
        RECT 296.200 139.475 296.370 140.415 ;
        RECT 296.640 139.475 296.810 141.125 ;
        RECT 297.480 139.475 297.650 140.415 ;
        RECT 298.180 139.535 298.570 141.125 ;
        RECT 298.940 139.475 299.110 141.125 ;
        RECT 299.380 139.475 299.550 140.415 ;
        RECT 299.820 139.475 299.990 141.125 ;
        RECT 300.160 139.475 300.430 140.415 ;
        RECT 300.700 139.475 300.870 141.125 ;
        RECT 301.585 139.475 301.755 141.125 ;
        RECT 302.025 139.475 302.195 140.415 ;
        RECT 302.465 139.475 302.635 141.125 ;
        RECT 303.180 139.535 303.570 141.125 ;
        RECT 304.085 139.475 304.255 141.125 ;
        RECT 304.525 139.475 304.695 140.415 ;
        RECT 304.965 139.475 305.135 141.125 ;
        RECT 305.835 139.475 306.005 141.125 ;
        RECT 306.275 139.475 306.445 140.415 ;
        RECT 306.715 139.475 306.885 141.125 ;
        RECT 307.585 139.475 307.755 141.125 ;
        RECT 308.025 139.475 308.195 140.415 ;
        RECT 308.465 139.475 308.635 141.125 ;
        RECT 309.335 139.475 309.505 141.125 ;
        RECT 309.775 139.475 309.945 140.415 ;
        RECT 310.215 139.475 310.385 141.125 ;
        RECT 310.930 139.535 311.320 141.125 ;
        RECT 316.030 140.630 316.750 140.800 ;
        RECT 316.030 139.770 316.200 140.630 ;
        RECT 294.365 139.185 295.220 139.265 ;
        RECT 294.365 138.855 295.250 139.185 ;
        RECT 296.280 139.005 296.620 139.260 ;
        RECT 297.420 139.090 297.750 139.305 ;
        RECT 299.430 139.095 300.120 139.265 ;
        RECT 299.430 139.050 299.760 139.095 ;
        RECT 300.460 139.090 301.000 139.305 ;
        RECT 301.865 139.185 302.720 139.265 ;
        RECT 304.365 139.185 305.220 139.265 ;
        RECT 306.115 139.185 306.970 139.265 ;
        RECT 307.865 139.185 308.720 139.265 ;
        RECT 309.615 139.185 310.470 139.265 ;
        RECT 299.940 138.905 300.270 138.925 ;
        RECT 294.365 138.775 295.220 138.855 ;
        RECT 296.760 138.735 297.690 138.905 ;
        RECT 299.940 138.735 300.940 138.905 ;
        RECT 301.865 138.855 302.750 139.185 ;
        RECT 304.365 138.855 305.250 139.185 ;
        RECT 306.115 138.855 307.000 139.185 ;
        RECT 307.865 138.855 308.750 139.185 ;
        RECT 309.615 138.855 310.500 139.185 ;
        RECT 301.865 138.775 302.720 138.855 ;
        RECT 304.365 138.775 305.220 138.855 ;
        RECT 306.115 138.775 306.970 138.855 ;
        RECT 307.865 138.775 308.720 138.855 ;
        RECT 309.615 138.775 310.470 138.855 ;
        RECT 293.180 137.365 293.570 138.730 ;
        RECT 294.085 137.365 294.255 138.565 ;
        RECT 294.525 138.075 294.695 138.565 ;
        RECT 294.965 137.365 295.135 138.565 ;
        RECT 295.760 137.365 295.930 138.565 ;
        RECT 296.200 138.075 296.370 138.565 ;
        RECT 296.640 137.365 296.810 138.565 ;
        RECT 297.080 137.910 297.250 138.565 ;
        RECT 297.520 137.365 297.690 138.565 ;
        RECT 298.180 137.365 298.570 138.730 ;
        RECT 298.940 137.365 299.110 138.565 ;
        RECT 299.380 138.075 299.550 138.565 ;
        RECT 299.820 137.365 299.990 138.565 ;
        RECT 300.160 138.075 300.830 138.565 ;
        RECT 301.585 137.365 301.755 138.565 ;
        RECT 302.025 138.075 302.195 138.565 ;
        RECT 302.465 137.365 302.635 138.565 ;
        RECT 303.180 137.365 303.570 138.730 ;
        RECT 304.085 137.365 304.255 138.565 ;
        RECT 304.525 138.075 304.695 138.565 ;
        RECT 304.965 137.365 305.135 138.565 ;
        RECT 305.835 137.365 306.005 138.565 ;
        RECT 306.275 138.075 306.445 138.565 ;
        RECT 306.715 137.365 306.885 138.565 ;
        RECT 307.585 137.365 307.755 138.565 ;
        RECT 308.025 138.075 308.195 138.565 ;
        RECT 308.465 137.365 308.635 138.565 ;
        RECT 309.335 137.365 309.505 138.565 ;
        RECT 309.775 138.075 309.945 138.565 ;
        RECT 310.215 137.365 310.385 138.565 ;
        RECT 310.930 137.365 311.320 138.730 ;
        RECT 315.660 137.640 315.830 139.730 ;
        RECT 316.000 138.735 316.170 139.065 ;
        RECT 316.370 138.920 316.540 140.415 ;
        RECT 316.870 139.260 317.040 140.460 ;
        RECT 317.210 139.475 317.380 141.125 ;
        RECT 317.550 140.660 317.880 140.955 ;
        RECT 317.650 139.260 317.820 140.415 ;
        RECT 318.090 139.475 318.260 141.125 ;
        RECT 318.430 140.630 318.760 140.800 ;
        RECT 318.530 139.475 318.920 140.415 ;
        RECT 319.090 139.475 319.260 141.125 ;
        RECT 319.530 139.475 319.700 140.415 ;
        RECT 319.970 139.475 320.140 141.125 ;
        RECT 320.680 139.535 321.070 141.125 ;
        RECT 321.615 139.475 321.785 141.125 ;
        RECT 322.055 139.475 322.225 140.415 ;
        RECT 322.495 139.475 322.665 141.125 ;
        RECT 323.485 139.475 323.655 141.125 ;
        RECT 323.925 139.475 324.195 140.415 ;
        RECT 324.365 139.475 324.535 141.125 ;
        RECT 324.705 140.660 325.035 140.955 ;
        RECT 325.445 140.785 325.775 140.955 ;
        RECT 325.525 140.660 325.695 140.785 ;
        RECT 324.805 139.475 324.975 140.460 ;
        RECT 316.870 139.090 317.480 139.260 ;
        RECT 317.650 139.090 318.080 139.260 ;
        RECT 316.370 138.750 317.700 138.920 ;
        RECT 316.010 138.075 316.180 138.565 ;
        RECT 316.450 137.365 316.620 138.565 ;
        RECT 316.790 138.315 316.960 138.750 ;
        RECT 317.910 138.565 318.080 139.090 ;
        RECT 317.210 138.155 317.540 138.485 ;
        RECT 317.850 138.075 318.080 138.565 ;
        RECT 318.250 137.905 318.420 138.920 ;
        RECT 318.750 138.905 318.920 139.475 ;
        RECT 319.130 139.090 319.680 139.260 ;
        RECT 321.530 139.185 322.385 139.265 ;
        RECT 318.750 138.735 319.140 138.905 ;
        RECT 321.500 138.855 322.385 139.185 ;
        RECT 323.310 139.135 323.850 139.305 ;
        RECT 321.530 138.775 322.385 138.855 ;
        RECT 323.670 138.735 323.850 139.135 ;
        RECT 318.750 138.315 318.920 138.735 ;
        RECT 316.790 137.535 317.120 137.840 ;
        RECT 317.940 137.735 318.420 137.905 ;
        RECT 318.590 137.535 318.920 137.840 ;
        RECT 319.090 137.365 319.260 138.565 ;
        RECT 319.530 138.075 319.700 138.565 ;
        RECT 319.970 137.365 320.140 138.565 ;
        RECT 320.680 137.365 321.070 138.730 ;
        RECT 324.020 138.565 324.195 139.475 ;
        RECT 324.365 138.935 325.075 139.305 ;
        RECT 321.615 137.365 321.785 138.565 ;
        RECT 322.055 138.075 322.225 138.565 ;
        RECT 322.495 137.365 322.665 138.565 ;
        RECT 323.525 137.365 323.695 138.565 ;
        RECT 323.965 138.075 324.195 138.565 ;
        RECT 324.405 137.365 324.575 138.565 ;
        RECT 324.905 137.705 325.075 138.210 ;
        RECT 325.245 138.075 325.515 140.415 ;
        RECT 325.685 139.475 325.855 140.460 ;
        RECT 326.125 139.475 326.295 141.125 ;
        RECT 325.875 138.735 326.355 139.260 ;
        RECT 324.745 137.535 325.075 137.705 ;
        RECT 325.365 137.670 325.695 137.905 ;
        RECT 326.085 137.365 326.255 138.565 ;
        RECT 326.525 138.075 326.795 140.415 ;
        RECT 327.005 139.475 327.175 141.125 ;
        RECT 327.680 139.535 328.070 141.125 ;
        RECT 329.030 140.630 329.750 140.800 ;
        RECT 329.030 139.770 329.200 140.630 ;
        RECT 326.965 137.365 327.135 138.565 ;
        RECT 327.680 137.365 328.070 138.730 ;
        RECT 328.660 137.640 328.830 139.730 ;
        RECT 329.000 138.735 329.170 139.065 ;
        RECT 329.370 138.920 329.540 140.415 ;
        RECT 329.870 139.260 330.040 140.460 ;
        RECT 330.210 139.475 330.380 141.125 ;
        RECT 330.550 140.660 330.880 140.955 ;
        RECT 330.650 139.260 330.820 140.415 ;
        RECT 331.090 139.475 331.260 141.125 ;
        RECT 331.430 140.630 331.760 140.800 ;
        RECT 331.530 139.475 331.920 140.415 ;
        RECT 332.090 139.475 332.260 141.125 ;
        RECT 332.530 139.475 332.700 140.415 ;
        RECT 332.970 139.475 333.140 141.125 ;
        RECT 333.680 139.535 334.070 141.125 ;
        RECT 334.615 139.475 334.785 141.125 ;
        RECT 335.055 139.475 335.225 140.415 ;
        RECT 335.495 139.475 335.665 141.125 ;
        RECT 336.485 139.475 336.655 141.125 ;
        RECT 336.925 139.475 337.195 140.415 ;
        RECT 337.365 139.475 337.535 141.125 ;
        RECT 337.705 140.660 338.035 140.955 ;
        RECT 338.445 140.785 338.775 140.955 ;
        RECT 338.525 140.660 338.695 140.785 ;
        RECT 337.805 139.475 337.975 140.460 ;
        RECT 329.870 139.090 330.480 139.260 ;
        RECT 330.650 139.090 331.080 139.260 ;
        RECT 329.370 138.750 330.700 138.920 ;
        RECT 329.010 138.075 329.180 138.565 ;
        RECT 329.450 137.365 329.620 138.565 ;
        RECT 329.790 138.315 329.960 138.750 ;
        RECT 330.910 138.565 331.080 139.090 ;
        RECT 330.210 138.155 330.540 138.485 ;
        RECT 330.850 138.075 331.080 138.565 ;
        RECT 331.250 137.905 331.420 138.920 ;
        RECT 331.750 138.905 331.920 139.475 ;
        RECT 332.130 139.090 332.680 139.260 ;
        RECT 334.530 139.185 335.385 139.265 ;
        RECT 331.750 138.735 332.140 138.905 ;
        RECT 334.500 138.855 335.385 139.185 ;
        RECT 336.310 139.135 336.850 139.305 ;
        RECT 334.530 138.775 335.385 138.855 ;
        RECT 336.670 138.735 336.850 139.135 ;
        RECT 331.750 138.315 331.920 138.735 ;
        RECT 329.790 137.535 330.120 137.840 ;
        RECT 330.940 137.735 331.420 137.905 ;
        RECT 331.590 137.535 331.920 137.840 ;
        RECT 332.090 137.365 332.260 138.565 ;
        RECT 332.530 138.075 332.700 138.565 ;
        RECT 332.970 137.365 333.140 138.565 ;
        RECT 333.680 137.365 334.070 138.730 ;
        RECT 337.020 138.565 337.195 139.475 ;
        RECT 337.365 138.935 338.075 139.305 ;
        RECT 334.615 137.365 334.785 138.565 ;
        RECT 335.055 138.075 335.225 138.565 ;
        RECT 335.495 137.365 335.665 138.565 ;
        RECT 336.525 137.365 336.695 138.565 ;
        RECT 336.965 138.075 337.195 138.565 ;
        RECT 337.405 137.365 337.575 138.565 ;
        RECT 337.905 137.705 338.075 138.210 ;
        RECT 338.245 138.075 338.515 140.415 ;
        RECT 338.685 139.475 338.855 140.460 ;
        RECT 339.125 139.475 339.295 141.125 ;
        RECT 338.875 138.735 339.355 139.260 ;
        RECT 337.745 137.535 338.075 137.705 ;
        RECT 338.365 137.670 338.695 137.905 ;
        RECT 339.085 137.365 339.255 138.565 ;
        RECT 339.525 138.075 339.795 140.415 ;
        RECT 340.005 139.475 340.175 141.125 ;
        RECT 340.680 139.535 341.070 141.125 ;
        RECT 343.990 139.475 344.160 141.125 ;
        RECT 344.430 139.475 344.600 140.415 ;
        RECT 344.870 139.475 345.040 141.125 ;
        RECT 345.615 139.475 345.785 141.125 ;
        RECT 346.055 139.475 346.225 140.415 ;
        RECT 346.495 139.475 346.665 141.125 ;
        RECT 347.115 139.475 347.285 141.125 ;
        RECT 347.555 139.475 347.725 140.415 ;
        RECT 347.995 139.475 348.165 141.125 ;
        RECT 348.680 139.535 349.070 141.125 ;
        RECT 349.615 139.475 349.785 141.125 ;
        RECT 350.055 139.475 350.225 140.415 ;
        RECT 350.495 139.475 350.665 141.125 ;
        RECT 343.815 139.075 344.880 139.305 ;
        RECT 345.530 139.185 346.385 139.265 ;
        RECT 347.030 139.185 347.885 139.265 ;
        RECT 349.530 139.185 350.385 139.265 ;
        RECT 343.810 138.735 344.400 138.905 ;
        RECT 345.500 138.855 346.385 139.185 ;
        RECT 347.000 138.855 347.885 139.185 ;
        RECT 349.500 138.855 350.385 139.185 ;
        RECT 345.530 138.775 346.385 138.855 ;
        RECT 347.030 138.775 347.885 138.855 ;
        RECT 349.530 138.775 350.385 138.855 ;
        RECT 339.965 137.365 340.135 138.565 ;
        RECT 340.680 137.365 341.070 138.730 ;
        RECT 343.990 137.365 344.160 138.565 ;
        RECT 344.830 138.075 345.000 138.565 ;
        RECT 345.615 137.365 345.785 138.565 ;
        RECT 346.055 138.075 346.225 138.565 ;
        RECT 346.495 137.365 346.665 138.565 ;
        RECT 347.115 137.365 347.285 138.565 ;
        RECT 347.555 138.075 347.725 138.565 ;
        RECT 347.995 137.365 348.165 138.565 ;
        RECT 348.680 137.365 349.070 138.730 ;
        RECT 349.615 137.365 349.785 138.565 ;
        RECT 350.055 138.075 350.225 138.565 ;
        RECT 350.495 137.365 350.665 138.565 ;
        RECT 293.000 137.115 341.250 137.365 ;
        RECT 343.500 137.115 351.000 137.365 ;
        RECT 292.750 134.125 351.000 134.375 ;
        RECT 292.930 132.535 293.320 134.125 ;
        RECT 293.860 132.475 294.030 134.125 ;
        RECT 294.300 132.475 294.470 133.415 ;
        RECT 294.740 132.475 294.910 134.125 ;
        RECT 295.240 133.630 295.570 133.800 ;
        RECT 295.080 132.475 295.470 133.415 ;
        RECT 295.740 132.475 295.910 134.125 ;
        RECT 296.120 133.660 296.450 133.955 ;
        RECT 294.320 132.090 294.870 132.260 ;
        RECT 295.080 131.905 295.250 132.475 ;
        RECT 296.180 132.260 296.350 133.415 ;
        RECT 296.620 132.475 296.790 134.125 ;
        RECT 297.250 133.630 297.970 133.800 ;
        RECT 296.960 132.260 297.130 133.460 ;
        RECT 295.920 132.090 296.350 132.260 ;
        RECT 296.520 132.090 297.130 132.260 ;
        RECT 294.860 131.735 295.250 131.905 ;
        RECT 292.930 130.365 293.320 131.730 ;
        RECT 293.860 130.365 294.030 131.565 ;
        RECT 294.300 131.075 294.470 131.565 ;
        RECT 294.740 130.365 294.910 131.565 ;
        RECT 295.080 131.315 295.250 131.735 ;
        RECT 295.580 130.905 295.750 131.920 ;
        RECT 295.920 131.565 296.090 132.090 ;
        RECT 297.460 131.920 297.630 133.415 ;
        RECT 297.800 132.770 297.970 133.630 ;
        RECT 296.300 131.750 297.630 131.920 ;
        RECT 295.920 131.075 296.150 131.565 ;
        RECT 296.460 131.155 296.790 131.485 ;
        RECT 297.040 131.315 297.210 131.750 ;
        RECT 297.830 131.735 298.000 132.065 ;
        RECT 295.080 130.535 295.410 130.840 ;
        RECT 295.580 130.735 296.060 130.905 ;
        RECT 296.880 130.535 297.210 130.840 ;
        RECT 297.380 130.365 297.550 131.565 ;
        RECT 297.820 131.075 297.990 131.565 ;
        RECT 298.170 130.640 298.340 132.730 ;
        RECT 298.940 132.475 299.110 134.125 ;
        RECT 299.380 132.475 299.550 133.415 ;
        RECT 299.820 132.475 299.990 134.125 ;
        RECT 300.160 132.475 300.430 133.415 ;
        RECT 300.700 132.475 300.870 134.125 ;
        RECT 301.585 132.475 301.755 134.125 ;
        RECT 302.025 132.475 302.195 133.415 ;
        RECT 302.465 132.475 302.635 134.125 ;
        RECT 303.180 132.535 303.570 134.125 ;
        RECT 304.085 132.475 304.255 134.125 ;
        RECT 304.525 132.475 304.695 133.415 ;
        RECT 304.965 132.475 305.135 134.125 ;
        RECT 305.835 132.475 306.005 134.125 ;
        RECT 306.275 132.475 306.445 133.415 ;
        RECT 306.715 132.475 306.885 134.125 ;
        RECT 307.585 132.475 307.755 134.125 ;
        RECT 308.025 132.475 308.195 133.415 ;
        RECT 308.465 132.475 308.635 134.125 ;
        RECT 309.335 132.475 309.505 134.125 ;
        RECT 309.775 132.475 309.945 133.415 ;
        RECT 310.215 132.475 310.385 134.125 ;
        RECT 310.930 132.535 311.320 134.125 ;
        RECT 311.770 132.475 311.940 134.125 ;
        RECT 312.210 132.475 312.380 133.415 ;
        RECT 312.650 132.475 312.820 134.125 ;
        RECT 313.030 133.660 313.360 133.955 ;
        RECT 313.090 132.305 313.260 133.415 ;
        RECT 313.530 132.475 313.700 134.125 ;
        RECT 313.870 133.660 314.200 133.955 ;
        RECT 313.970 132.305 314.140 133.415 ;
        RECT 314.410 132.475 314.580 134.125 ;
        RECT 299.430 132.095 300.120 132.265 ;
        RECT 299.430 132.050 299.760 132.095 ;
        RECT 300.460 132.090 301.000 132.305 ;
        RECT 301.865 132.185 302.720 132.265 ;
        RECT 304.365 132.185 305.220 132.265 ;
        RECT 306.115 132.185 306.970 132.265 ;
        RECT 307.865 132.185 308.720 132.265 ;
        RECT 309.615 132.185 310.470 132.265 ;
        RECT 299.940 131.905 300.270 131.925 ;
        RECT 299.940 131.735 300.940 131.905 ;
        RECT 301.865 131.855 302.750 132.185 ;
        RECT 304.365 131.855 305.250 132.185 ;
        RECT 306.115 131.855 307.000 132.185 ;
        RECT 307.865 131.855 308.750 132.185 ;
        RECT 309.615 131.855 310.500 132.185 ;
        RECT 312.000 132.135 314.140 132.305 ;
        RECT 312.000 132.090 312.620 132.135 ;
        RECT 312.770 131.905 313.100 131.965 ;
        RECT 301.865 131.775 302.720 131.855 ;
        RECT 304.365 131.775 305.220 131.855 ;
        RECT 306.115 131.775 306.970 131.855 ;
        RECT 307.865 131.775 308.720 131.855 ;
        RECT 309.615 131.775 310.470 131.855 ;
        RECT 312.770 131.735 313.580 131.905 ;
        RECT 314.010 131.795 314.340 131.965 ;
        RECT 298.940 130.365 299.110 131.565 ;
        RECT 299.380 131.075 299.550 131.565 ;
        RECT 299.820 130.365 299.990 131.565 ;
        RECT 300.160 131.075 300.830 131.565 ;
        RECT 301.585 130.365 301.755 131.565 ;
        RECT 302.025 131.075 302.195 131.565 ;
        RECT 302.465 130.365 302.635 131.565 ;
        RECT 303.180 130.365 303.570 131.730 ;
        RECT 304.085 130.365 304.255 131.565 ;
        RECT 304.525 131.075 304.695 131.565 ;
        RECT 304.965 130.365 305.135 131.565 ;
        RECT 305.835 130.365 306.005 131.565 ;
        RECT 306.275 131.075 306.445 131.565 ;
        RECT 306.715 130.365 306.885 131.565 ;
        RECT 307.585 130.365 307.755 131.565 ;
        RECT 308.025 131.075 308.195 131.565 ;
        RECT 308.465 130.365 308.635 131.565 ;
        RECT 309.335 130.365 309.505 131.565 ;
        RECT 309.775 131.075 309.945 131.565 ;
        RECT 310.215 130.365 310.385 131.565 ;
        RECT 310.930 130.365 311.320 131.730 ;
        RECT 311.770 130.365 311.940 131.565 ;
        RECT 312.210 131.075 312.380 131.565 ;
        RECT 312.650 130.365 312.820 131.565 ;
        RECT 313.010 130.705 313.180 131.565 ;
        RECT 313.410 131.270 313.580 131.735 ;
        RECT 314.290 131.045 314.460 131.565 ;
        RECT 313.600 130.875 314.460 131.045 ;
        RECT 314.750 130.705 314.920 133.480 ;
        RECT 315.430 132.535 315.820 134.125 ;
        RECT 316.325 132.475 316.495 134.125 ;
        RECT 313.010 130.535 313.430 130.705 ;
        RECT 313.680 130.535 314.920 130.705 ;
        RECT 315.430 130.365 315.820 131.730 ;
        RECT 316.365 130.365 316.535 131.565 ;
        RECT 316.705 131.075 316.975 133.415 ;
        RECT 317.205 132.475 317.375 134.125 ;
        RECT 317.725 133.785 318.055 133.955 ;
        RECT 317.805 133.660 317.975 133.785 ;
        RECT 318.465 133.660 318.795 133.955 ;
        RECT 317.645 132.475 317.815 133.460 ;
        RECT 317.145 131.735 317.625 132.260 ;
        RECT 317.245 130.365 317.415 131.565 ;
        RECT 317.985 131.075 318.255 133.415 ;
        RECT 318.525 132.475 318.695 133.460 ;
        RECT 318.965 132.475 319.135 134.125 ;
        RECT 319.305 132.475 319.575 133.415 ;
        RECT 319.845 132.475 320.015 134.125 ;
        RECT 320.835 132.475 321.005 134.125 ;
        RECT 321.275 132.475 321.445 133.415 ;
        RECT 321.715 132.475 321.885 134.125 ;
        RECT 322.430 132.535 322.820 134.125 ;
        RECT 323.360 132.475 323.530 134.125 ;
        RECT 323.800 132.475 323.970 133.415 ;
        RECT 324.240 132.475 324.410 134.125 ;
        RECT 324.740 133.630 325.070 133.800 ;
        RECT 324.580 132.475 324.970 133.415 ;
        RECT 325.240 132.475 325.410 134.125 ;
        RECT 325.620 133.660 325.950 133.955 ;
        RECT 318.425 131.935 319.135 132.305 ;
        RECT 319.305 131.565 319.480 132.475 ;
        RECT 319.650 132.135 320.190 132.305 ;
        RECT 321.115 132.185 321.970 132.265 ;
        RECT 319.650 131.735 319.830 132.135 ;
        RECT 321.115 131.855 322.000 132.185 ;
        RECT 323.820 132.090 324.370 132.260 ;
        RECT 324.580 131.905 324.750 132.475 ;
        RECT 325.680 132.260 325.850 133.415 ;
        RECT 326.120 132.475 326.290 134.125 ;
        RECT 326.750 133.630 327.470 133.800 ;
        RECT 326.460 132.260 326.630 133.460 ;
        RECT 325.420 132.090 325.850 132.260 ;
        RECT 326.020 132.090 326.630 132.260 ;
        RECT 321.115 131.775 321.970 131.855 ;
        RECT 324.360 131.735 324.750 131.905 ;
        RECT 317.805 130.670 318.135 130.905 ;
        RECT 318.425 130.705 318.595 131.210 ;
        RECT 318.425 130.535 318.755 130.705 ;
        RECT 318.925 130.365 319.095 131.565 ;
        RECT 319.305 131.075 319.535 131.565 ;
        RECT 319.805 130.365 319.975 131.565 ;
        RECT 320.835 130.365 321.005 131.565 ;
        RECT 321.275 131.075 321.445 131.565 ;
        RECT 321.715 130.365 321.885 131.565 ;
        RECT 322.430 130.365 322.820 131.730 ;
        RECT 323.360 130.365 323.530 131.565 ;
        RECT 323.800 131.075 323.970 131.565 ;
        RECT 324.240 130.365 324.410 131.565 ;
        RECT 324.580 131.315 324.750 131.735 ;
        RECT 325.080 130.905 325.250 131.920 ;
        RECT 325.420 131.565 325.590 132.090 ;
        RECT 326.960 131.920 327.130 133.415 ;
        RECT 327.300 132.770 327.470 133.630 ;
        RECT 325.800 131.750 327.130 131.920 ;
        RECT 325.420 131.075 325.650 131.565 ;
        RECT 325.960 131.155 326.290 131.485 ;
        RECT 326.540 131.315 326.710 131.750 ;
        RECT 327.330 131.735 327.500 132.065 ;
        RECT 324.580 130.535 324.910 130.840 ;
        RECT 325.080 130.735 325.560 130.905 ;
        RECT 326.380 130.535 326.710 130.840 ;
        RECT 326.880 130.365 327.050 131.565 ;
        RECT 327.320 131.075 327.490 131.565 ;
        RECT 327.670 130.640 327.840 132.730 ;
        RECT 328.430 132.535 328.820 134.125 ;
        RECT 329.325 132.475 329.495 134.125 ;
        RECT 328.430 130.365 328.820 131.730 ;
        RECT 329.365 130.365 329.535 131.565 ;
        RECT 329.705 131.075 329.975 133.415 ;
        RECT 330.205 132.475 330.375 134.125 ;
        RECT 330.725 133.785 331.055 133.955 ;
        RECT 330.805 133.660 330.975 133.785 ;
        RECT 331.465 133.660 331.795 133.955 ;
        RECT 330.645 132.475 330.815 133.460 ;
        RECT 330.145 131.735 330.625 132.260 ;
        RECT 330.245 130.365 330.415 131.565 ;
        RECT 330.985 131.075 331.255 133.415 ;
        RECT 331.525 132.475 331.695 133.460 ;
        RECT 331.965 132.475 332.135 134.125 ;
        RECT 332.305 132.475 332.575 133.415 ;
        RECT 332.845 132.475 333.015 134.125 ;
        RECT 333.835 132.475 334.005 134.125 ;
        RECT 334.275 132.475 334.445 133.415 ;
        RECT 334.715 132.475 334.885 134.125 ;
        RECT 335.430 132.535 335.820 134.125 ;
        RECT 336.360 132.475 336.530 134.125 ;
        RECT 336.800 132.475 336.970 133.415 ;
        RECT 337.240 132.475 337.410 134.125 ;
        RECT 337.740 133.630 338.070 133.800 ;
        RECT 337.580 132.475 337.970 133.415 ;
        RECT 338.240 132.475 338.410 134.125 ;
        RECT 338.620 133.660 338.950 133.955 ;
        RECT 331.425 131.935 332.135 132.305 ;
        RECT 332.305 131.565 332.480 132.475 ;
        RECT 332.650 132.135 333.190 132.305 ;
        RECT 334.115 132.185 334.970 132.265 ;
        RECT 332.650 131.735 332.830 132.135 ;
        RECT 334.115 131.855 335.000 132.185 ;
        RECT 336.820 132.090 337.370 132.260 ;
        RECT 337.580 131.905 337.750 132.475 ;
        RECT 338.680 132.260 338.850 133.415 ;
        RECT 339.120 132.475 339.290 134.125 ;
        RECT 339.750 133.630 340.470 133.800 ;
        RECT 339.460 132.260 339.630 133.460 ;
        RECT 338.420 132.090 338.850 132.260 ;
        RECT 339.020 132.090 339.630 132.260 ;
        RECT 334.115 131.775 334.970 131.855 ;
        RECT 337.360 131.735 337.750 131.905 ;
        RECT 330.805 130.670 331.135 130.905 ;
        RECT 331.425 130.705 331.595 131.210 ;
        RECT 331.425 130.535 331.755 130.705 ;
        RECT 331.925 130.365 332.095 131.565 ;
        RECT 332.305 131.075 332.535 131.565 ;
        RECT 332.805 130.365 332.975 131.565 ;
        RECT 333.835 130.365 334.005 131.565 ;
        RECT 334.275 131.075 334.445 131.565 ;
        RECT 334.715 130.365 334.885 131.565 ;
        RECT 335.430 130.365 335.820 131.730 ;
        RECT 336.360 130.365 336.530 131.565 ;
        RECT 336.800 131.075 336.970 131.565 ;
        RECT 337.240 130.365 337.410 131.565 ;
        RECT 337.580 131.315 337.750 131.735 ;
        RECT 338.080 130.905 338.250 131.920 ;
        RECT 338.420 131.565 338.590 132.090 ;
        RECT 339.960 131.920 340.130 133.415 ;
        RECT 340.300 132.770 340.470 133.630 ;
        RECT 338.800 131.750 340.130 131.920 ;
        RECT 338.420 131.075 338.650 131.565 ;
        RECT 338.960 131.155 339.290 131.485 ;
        RECT 339.540 131.315 339.710 131.750 ;
        RECT 340.330 131.735 340.500 132.065 ;
        RECT 337.580 130.535 337.910 130.840 ;
        RECT 338.080 130.735 338.560 130.905 ;
        RECT 339.380 130.535 339.710 130.840 ;
        RECT 339.880 130.365 340.050 131.565 ;
        RECT 340.320 131.075 340.490 131.565 ;
        RECT 340.670 130.640 340.840 132.730 ;
        RECT 341.430 132.535 341.820 134.125 ;
        RECT 342.365 132.475 342.535 134.125 ;
        RECT 342.805 132.475 342.975 133.415 ;
        RECT 343.245 132.475 343.415 134.125 ;
        RECT 343.990 132.475 344.160 134.125 ;
        RECT 344.430 132.475 344.600 133.415 ;
        RECT 344.870 132.475 345.040 134.125 ;
        RECT 345.615 132.475 345.785 134.125 ;
        RECT 346.055 132.475 346.225 133.415 ;
        RECT 346.495 132.475 346.665 134.125 ;
        RECT 347.115 132.475 347.285 134.125 ;
        RECT 347.555 132.475 347.725 133.415 ;
        RECT 347.995 132.475 348.165 134.125 ;
        RECT 348.680 132.535 349.070 134.125 ;
        RECT 349.615 132.475 349.785 134.125 ;
        RECT 350.055 132.475 350.225 133.415 ;
        RECT 350.495 132.475 350.665 134.125 ;
        RECT 342.280 132.185 343.135 132.265 ;
        RECT 342.250 131.855 343.135 132.185 ;
        RECT 343.815 132.075 344.880 132.305 ;
        RECT 345.530 132.185 346.385 132.265 ;
        RECT 347.030 132.185 347.885 132.265 ;
        RECT 349.530 132.185 350.385 132.265 ;
        RECT 342.280 131.775 343.135 131.855 ;
        RECT 343.810 131.735 344.400 131.905 ;
        RECT 345.500 131.855 346.385 132.185 ;
        RECT 347.000 131.855 347.885 132.185 ;
        RECT 349.500 131.855 350.385 132.185 ;
        RECT 345.530 131.775 346.385 131.855 ;
        RECT 347.030 131.775 347.885 131.855 ;
        RECT 349.530 131.775 350.385 131.855 ;
        RECT 341.430 130.365 341.820 131.730 ;
        RECT 342.365 130.365 342.535 131.565 ;
        RECT 342.805 131.075 342.975 131.565 ;
        RECT 343.245 130.365 343.415 131.565 ;
        RECT 343.990 130.365 344.160 131.565 ;
        RECT 344.830 131.075 345.000 131.565 ;
        RECT 345.615 130.365 345.785 131.565 ;
        RECT 346.055 131.075 346.225 131.565 ;
        RECT 346.495 130.365 346.665 131.565 ;
        RECT 347.115 130.365 347.285 131.565 ;
        RECT 347.555 131.075 347.725 131.565 ;
        RECT 347.995 130.365 348.165 131.565 ;
        RECT 348.680 130.365 349.070 131.730 ;
        RECT 349.615 130.365 349.785 131.565 ;
        RECT 350.055 131.075 350.225 131.565 ;
        RECT 350.495 130.365 350.665 131.565 ;
        RECT 292.750 130.115 351.000 130.365 ;
        RECT 354.000 127.250 354.500 151.250 ;
        RECT 390.875 151.375 391.125 157.625 ;
        RECT 393.915 156.750 394.085 157.250 ;
        RECT 391.615 151.730 391.785 155.770 ;
        RECT 392.075 151.730 392.245 155.770 ;
        RECT 392.535 151.730 392.705 155.770 ;
        RECT 392.995 151.730 393.165 155.770 ;
        RECT 393.455 151.730 393.625 155.770 ;
        RECT 393.915 151.730 394.085 155.770 ;
        RECT 394.375 151.730 394.545 155.770 ;
        RECT 394.835 151.730 395.005 155.770 ;
        RECT 395.295 151.730 395.465 155.770 ;
        RECT 395.755 151.730 395.925 155.770 ;
        RECT 396.215 151.730 396.385 155.770 ;
        RECT 396.875 151.375 397.125 157.625 ;
        RECT 399.915 156.750 400.085 157.250 ;
        RECT 397.615 151.730 397.785 155.770 ;
        RECT 398.075 151.730 398.245 155.770 ;
        RECT 398.535 151.730 398.705 155.770 ;
        RECT 398.995 151.730 399.165 155.770 ;
        RECT 399.455 151.730 399.625 155.770 ;
        RECT 399.915 151.730 400.085 155.770 ;
        RECT 400.375 151.730 400.545 155.770 ;
        RECT 400.835 151.730 401.005 155.770 ;
        RECT 401.295 151.730 401.465 155.770 ;
        RECT 401.755 151.730 401.925 155.770 ;
        RECT 402.215 151.730 402.385 155.770 ;
        RECT 402.875 151.375 403.125 157.625 ;
        RECT 405.915 156.750 406.085 157.250 ;
        RECT 403.615 151.730 403.785 155.770 ;
        RECT 404.075 151.730 404.245 155.770 ;
        RECT 404.535 151.730 404.705 155.770 ;
        RECT 404.995 151.730 405.165 155.770 ;
        RECT 405.455 151.730 405.625 155.770 ;
        RECT 405.915 151.730 406.085 155.770 ;
        RECT 406.375 151.730 406.545 155.770 ;
        RECT 406.835 151.730 407.005 155.770 ;
        RECT 407.295 151.730 407.465 155.770 ;
        RECT 407.755 151.730 407.925 155.770 ;
        RECT 408.215 151.730 408.385 155.770 ;
        RECT 408.875 151.375 409.125 157.625 ;
        RECT 409.625 157.625 420.875 157.875 ;
        RECT 409.625 153.375 409.875 157.625 ;
        RECT 412.415 156.750 412.585 157.250 ;
        RECT 410.215 153.805 410.385 155.845 ;
        RECT 410.655 153.805 410.825 155.845 ;
        RECT 411.095 153.805 411.265 155.845 ;
        RECT 411.535 153.805 411.705 155.845 ;
        RECT 411.975 153.805 412.145 155.845 ;
        RECT 412.415 153.805 412.585 155.845 ;
        RECT 412.855 153.805 413.025 155.845 ;
        RECT 413.295 153.805 413.465 155.845 ;
        RECT 413.735 153.805 413.905 155.845 ;
        RECT 414.175 153.805 414.345 155.845 ;
        RECT 414.615 153.805 414.785 155.845 ;
        RECT 415.125 153.375 415.375 157.625 ;
        RECT 417.915 156.750 418.085 157.250 ;
        RECT 415.715 153.805 415.885 155.845 ;
        RECT 416.155 153.805 416.325 155.845 ;
        RECT 416.595 153.805 416.765 155.845 ;
        RECT 417.035 153.805 417.205 155.845 ;
        RECT 417.475 153.805 417.645 155.845 ;
        RECT 417.915 153.805 418.085 155.845 ;
        RECT 418.355 153.805 418.525 155.845 ;
        RECT 418.795 153.805 418.965 155.845 ;
        RECT 419.235 153.805 419.405 155.845 ;
        RECT 419.675 153.805 419.845 155.845 ;
        RECT 420.115 153.805 420.285 155.845 ;
        RECT 420.625 153.375 420.875 157.625 ;
        RECT 409.625 153.125 420.875 153.375 ;
        RECT 390.875 151.125 409.125 151.375 ;
        RECT 286.250 126.750 354.500 127.250 ;
        RECT 388.125 149.875 391.375 150.125 ;
        RECT 388.125 146.375 388.375 149.875 ;
        RECT 389.665 149.000 389.835 149.500 ;
        RECT 388.780 147.730 389.260 148.770 ;
        RECT 389.530 147.730 389.970 148.770 ;
        RECT 390.240 147.730 390.720 148.770 ;
        RECT 389.665 147.000 389.835 147.500 ;
        RECT 391.125 146.375 391.375 149.875 ;
        RECT 388.125 146.125 391.375 146.375 ;
        RECT 388.125 142.625 388.375 146.125 ;
        RECT 389.665 145.250 389.835 145.750 ;
        RECT 388.780 143.980 389.260 145.020 ;
        RECT 389.530 143.980 389.970 145.020 ;
        RECT 390.240 143.980 390.720 145.020 ;
        RECT 389.665 143.250 389.835 143.750 ;
        RECT 391.125 142.625 391.375 146.125 ;
        RECT 388.125 142.375 391.375 142.625 ;
        RECT 388.125 138.875 388.375 142.375 ;
        RECT 389.665 141.500 389.835 142.000 ;
        RECT 388.780 140.230 389.260 141.270 ;
        RECT 389.530 140.230 389.970 141.270 ;
        RECT 390.240 140.230 390.720 141.270 ;
        RECT 389.665 139.500 389.835 140.000 ;
        RECT 391.125 138.875 391.375 142.375 ;
        RECT 388.125 138.625 391.375 138.875 ;
        RECT 388.125 135.125 388.375 138.625 ;
        RECT 389.665 137.750 389.835 138.250 ;
        RECT 388.780 136.480 389.260 137.520 ;
        RECT 389.530 136.480 389.970 137.520 ;
        RECT 390.240 136.480 390.720 137.520 ;
        RECT 389.665 135.750 389.835 136.250 ;
        RECT 391.125 135.125 391.375 138.625 ;
        RECT 388.125 134.875 391.375 135.125 ;
        RECT 388.125 131.375 388.375 134.875 ;
        RECT 389.665 134.000 389.835 134.500 ;
        RECT 388.780 132.730 389.260 133.770 ;
        RECT 389.530 132.730 389.970 133.770 ;
        RECT 390.240 132.730 390.720 133.770 ;
        RECT 389.665 132.000 389.835 132.500 ;
        RECT 391.125 131.375 391.375 134.875 ;
        RECT 388.125 131.125 391.375 131.375 ;
        RECT 388.125 127.625 388.375 131.125 ;
        RECT 389.665 130.250 389.835 130.750 ;
        RECT 388.780 128.980 389.260 130.020 ;
        RECT 389.530 128.980 389.970 130.020 ;
        RECT 390.240 128.980 390.720 130.020 ;
        RECT 389.665 128.250 389.835 128.750 ;
        RECT 391.125 127.625 391.375 131.125 ;
        RECT 388.125 127.375 391.375 127.625 ;
        RECT 294.250 125.750 350.250 126.250 ;
        RECT 294.250 112.750 294.750 125.750 ;
        RECT 298.500 123.875 346.500 124.125 ;
        RECT 298.780 122.750 298.950 123.580 ;
        RECT 299.320 123.380 299.650 123.550 ;
        RECT 298.780 122.250 299.070 122.750 ;
        RECT 298.780 120.435 298.950 122.250 ;
        RECT 299.240 122.225 299.630 123.165 ;
        RECT 300.080 122.225 300.250 123.875 ;
        RECT 300.580 123.380 300.910 123.550 ;
        RECT 300.640 122.225 300.910 123.165 ;
        RECT 301.080 122.225 301.250 123.875 ;
        RECT 299.120 121.605 299.290 121.935 ;
        RECT 299.460 121.855 299.630 122.225 ;
        RECT 300.740 121.935 300.910 122.225 ;
        RECT 301.520 121.935 301.690 123.165 ;
        RECT 302.080 122.225 302.250 123.875 ;
        RECT 302.520 122.225 302.790 123.165 ;
        RECT 302.960 122.225 303.130 123.875 ;
        RECT 303.865 122.225 304.035 123.875 ;
        RECT 304.305 122.225 304.475 123.165 ;
        RECT 304.745 122.225 304.915 123.875 ;
        RECT 305.600 122.225 305.770 123.875 ;
        RECT 306.440 122.225 306.610 123.165 ;
        RECT 307.180 122.285 307.570 123.875 ;
        RECT 308.100 122.225 308.270 123.875 ;
        RECT 308.940 122.225 309.110 123.165 ;
        RECT 309.780 122.750 309.950 123.580 ;
        RECT 310.320 123.380 310.650 123.550 ;
        RECT 309.780 122.250 310.070 122.750 ;
        RECT 299.460 121.685 300.570 121.855 ;
        RECT 299.460 121.315 299.630 121.685 ;
        RECT 300.740 121.610 301.350 121.935 ;
        RECT 300.740 121.315 300.910 121.610 ;
        RECT 301.180 121.605 301.350 121.610 ;
        RECT 301.520 121.605 302.450 121.935 ;
        RECT 301.520 121.315 301.690 121.605 ;
        RECT 302.620 121.315 302.790 122.225 ;
        RECT 303.780 121.935 304.635 122.015 ;
        RECT 303.750 121.605 304.635 121.935 ;
        RECT 305.500 121.840 305.830 122.055 ;
        RECT 306.000 121.885 306.690 122.055 ;
        RECT 303.780 121.525 304.635 121.605 ;
        RECT 299.360 120.825 299.630 121.315 ;
        RECT 299.800 120.115 299.970 121.315 ;
        RECT 300.640 120.825 300.910 121.315 ;
        RECT 301.240 121.145 301.690 121.315 ;
        RECT 301.240 120.825 301.410 121.145 ;
        RECT 300.140 120.285 301.650 120.635 ;
        RECT 302.080 120.115 302.250 121.315 ;
        RECT 302.520 120.825 302.790 121.315 ;
        RECT 302.960 120.115 303.130 121.315 ;
        RECT 303.865 120.115 304.035 121.315 ;
        RECT 304.305 120.825 304.475 121.315 ;
        RECT 304.745 120.115 304.915 121.315 ;
        RECT 305.560 120.115 305.730 121.315 ;
        RECT 306.000 120.825 306.170 121.885 ;
        RECT 308.000 121.840 308.330 122.055 ;
        RECT 308.500 121.885 309.190 122.055 ;
        RECT 306.340 121.485 306.670 121.655 ;
        RECT 306.440 120.115 306.610 121.315 ;
        RECT 307.180 120.115 307.570 121.480 ;
        RECT 308.060 120.115 308.230 121.315 ;
        RECT 308.500 120.825 308.670 121.885 ;
        RECT 308.840 121.485 309.170 121.655 ;
        RECT 308.940 120.115 309.110 121.315 ;
        RECT 309.780 120.435 309.950 122.250 ;
        RECT 310.240 122.225 310.630 123.165 ;
        RECT 311.080 122.225 311.250 123.875 ;
        RECT 311.580 123.380 311.910 123.550 ;
        RECT 311.640 122.225 311.910 123.165 ;
        RECT 312.080 122.225 312.250 123.875 ;
        RECT 310.120 121.605 310.290 121.935 ;
        RECT 310.460 121.855 310.630 122.225 ;
        RECT 311.740 121.935 311.910 122.225 ;
        RECT 312.520 121.935 312.690 123.165 ;
        RECT 313.080 122.225 313.250 123.875 ;
        RECT 313.520 122.225 313.790 123.165 ;
        RECT 313.960 122.225 314.130 123.875 ;
        RECT 314.780 122.750 314.950 123.580 ;
        RECT 315.320 123.380 315.650 123.550 ;
        RECT 314.780 122.250 315.070 122.750 ;
        RECT 310.460 121.685 311.570 121.855 ;
        RECT 310.460 121.315 310.630 121.685 ;
        RECT 311.740 121.610 312.350 121.935 ;
        RECT 311.740 121.315 311.910 121.610 ;
        RECT 312.180 121.605 312.350 121.610 ;
        RECT 312.520 121.605 313.450 121.935 ;
        RECT 312.520 121.315 312.690 121.605 ;
        RECT 313.620 121.315 313.790 122.225 ;
        RECT 310.360 120.825 310.630 121.315 ;
        RECT 310.800 120.115 310.970 121.315 ;
        RECT 311.640 120.825 311.910 121.315 ;
        RECT 312.240 121.145 312.690 121.315 ;
        RECT 312.240 120.825 312.410 121.145 ;
        RECT 311.140 120.285 312.650 120.635 ;
        RECT 313.080 120.115 313.250 121.315 ;
        RECT 313.520 120.825 313.790 121.315 ;
        RECT 313.960 120.115 314.130 121.315 ;
        RECT 314.780 120.435 314.950 122.250 ;
        RECT 315.240 122.225 315.630 123.165 ;
        RECT 316.080 122.225 316.250 123.875 ;
        RECT 316.580 123.380 316.910 123.550 ;
        RECT 316.640 122.225 316.910 123.165 ;
        RECT 317.080 122.225 317.250 123.875 ;
        RECT 315.120 121.605 315.290 121.935 ;
        RECT 315.460 121.855 315.630 122.225 ;
        RECT 316.740 121.935 316.910 122.225 ;
        RECT 317.520 121.935 317.690 123.165 ;
        RECT 318.080 122.225 318.250 123.875 ;
        RECT 318.520 122.225 318.790 123.165 ;
        RECT 318.960 122.225 319.130 123.875 ;
        RECT 319.865 122.225 320.035 123.875 ;
        RECT 320.305 122.225 320.475 123.165 ;
        RECT 320.745 122.225 320.915 123.875 ;
        RECT 321.600 122.225 321.770 123.875 ;
        RECT 322.440 122.225 322.610 123.165 ;
        RECT 323.180 122.285 323.570 123.875 ;
        RECT 324.100 122.225 324.270 123.875 ;
        RECT 324.940 122.225 325.110 123.165 ;
        RECT 325.780 122.750 325.950 123.580 ;
        RECT 326.320 123.380 326.650 123.550 ;
        RECT 325.780 122.250 326.070 122.750 ;
        RECT 315.460 121.685 316.570 121.855 ;
        RECT 315.460 121.315 315.630 121.685 ;
        RECT 316.740 121.610 317.350 121.935 ;
        RECT 316.740 121.315 316.910 121.610 ;
        RECT 317.180 121.605 317.350 121.610 ;
        RECT 317.520 121.605 318.450 121.935 ;
        RECT 317.520 121.315 317.690 121.605 ;
        RECT 318.620 121.315 318.790 122.225 ;
        RECT 319.780 121.935 320.635 122.015 ;
        RECT 319.750 121.605 320.635 121.935 ;
        RECT 321.500 121.840 321.830 122.055 ;
        RECT 322.000 121.885 322.690 122.055 ;
        RECT 319.780 121.525 320.635 121.605 ;
        RECT 315.360 120.825 315.630 121.315 ;
        RECT 315.800 120.115 315.970 121.315 ;
        RECT 316.640 120.825 316.910 121.315 ;
        RECT 317.240 121.145 317.690 121.315 ;
        RECT 317.240 120.825 317.410 121.145 ;
        RECT 316.140 120.285 317.650 120.635 ;
        RECT 318.080 120.115 318.250 121.315 ;
        RECT 318.520 120.825 318.790 121.315 ;
        RECT 318.960 120.115 319.130 121.315 ;
        RECT 319.865 120.115 320.035 121.315 ;
        RECT 320.305 120.825 320.475 121.315 ;
        RECT 320.745 120.115 320.915 121.315 ;
        RECT 321.560 120.115 321.730 121.315 ;
        RECT 322.000 120.825 322.170 121.885 ;
        RECT 324.000 121.840 324.330 122.055 ;
        RECT 324.500 121.885 325.190 122.055 ;
        RECT 322.340 121.485 322.670 121.655 ;
        RECT 322.440 120.115 322.610 121.315 ;
        RECT 323.180 120.115 323.570 121.480 ;
        RECT 324.060 120.115 324.230 121.315 ;
        RECT 324.500 120.825 324.670 121.885 ;
        RECT 324.840 121.485 325.170 121.655 ;
        RECT 324.940 120.115 325.110 121.315 ;
        RECT 325.780 120.435 325.950 122.250 ;
        RECT 326.240 122.225 326.630 123.165 ;
        RECT 327.080 122.225 327.250 123.875 ;
        RECT 327.580 123.380 327.910 123.550 ;
        RECT 327.640 122.225 327.910 123.165 ;
        RECT 328.080 122.225 328.250 123.875 ;
        RECT 326.120 121.605 326.290 121.935 ;
        RECT 326.460 121.855 326.630 122.225 ;
        RECT 327.740 121.935 327.910 122.225 ;
        RECT 328.520 121.935 328.690 123.165 ;
        RECT 329.080 122.225 329.250 123.875 ;
        RECT 329.520 122.225 329.790 123.165 ;
        RECT 329.960 122.225 330.130 123.875 ;
        RECT 330.780 122.750 330.950 123.580 ;
        RECT 331.320 123.380 331.650 123.550 ;
        RECT 330.780 122.250 331.070 122.750 ;
        RECT 326.460 121.685 327.570 121.855 ;
        RECT 326.460 121.315 326.630 121.685 ;
        RECT 327.740 121.610 328.350 121.935 ;
        RECT 327.740 121.315 327.910 121.610 ;
        RECT 328.180 121.605 328.350 121.610 ;
        RECT 328.520 121.605 329.450 121.935 ;
        RECT 328.520 121.315 328.690 121.605 ;
        RECT 329.620 121.315 329.790 122.225 ;
        RECT 326.360 120.825 326.630 121.315 ;
        RECT 326.800 120.115 326.970 121.315 ;
        RECT 327.640 120.825 327.910 121.315 ;
        RECT 328.240 121.145 328.690 121.315 ;
        RECT 328.240 120.825 328.410 121.145 ;
        RECT 327.140 120.285 328.650 120.635 ;
        RECT 329.080 120.115 329.250 121.315 ;
        RECT 329.520 120.825 329.790 121.315 ;
        RECT 329.960 120.115 330.130 121.315 ;
        RECT 330.780 120.435 330.950 122.250 ;
        RECT 331.240 122.225 331.630 123.165 ;
        RECT 332.080 122.225 332.250 123.875 ;
        RECT 332.580 123.380 332.910 123.550 ;
        RECT 332.640 122.225 332.910 123.165 ;
        RECT 333.080 122.225 333.250 123.875 ;
        RECT 331.120 121.605 331.290 121.935 ;
        RECT 331.460 121.855 331.630 122.225 ;
        RECT 332.740 121.935 332.910 122.225 ;
        RECT 333.520 121.935 333.690 123.165 ;
        RECT 334.080 122.225 334.250 123.875 ;
        RECT 334.520 122.225 334.790 123.165 ;
        RECT 334.960 122.225 335.130 123.875 ;
        RECT 335.865 122.225 336.035 123.875 ;
        RECT 336.305 122.225 336.475 123.165 ;
        RECT 336.745 122.225 336.915 123.875 ;
        RECT 337.600 122.225 337.770 123.875 ;
        RECT 338.440 122.225 338.610 123.165 ;
        RECT 339.180 122.285 339.570 123.875 ;
        RECT 340.100 122.225 340.270 123.875 ;
        RECT 340.940 122.225 341.110 123.165 ;
        RECT 341.780 122.750 341.950 123.580 ;
        RECT 342.320 123.380 342.650 123.550 ;
        RECT 341.780 122.250 342.070 122.750 ;
        RECT 331.460 121.685 332.570 121.855 ;
        RECT 331.460 121.315 331.630 121.685 ;
        RECT 332.740 121.610 333.350 121.935 ;
        RECT 332.740 121.315 332.910 121.610 ;
        RECT 333.180 121.605 333.350 121.610 ;
        RECT 333.520 121.605 334.450 121.935 ;
        RECT 333.520 121.315 333.690 121.605 ;
        RECT 334.620 121.315 334.790 122.225 ;
        RECT 335.780 121.935 336.635 122.015 ;
        RECT 335.750 121.605 336.635 121.935 ;
        RECT 337.500 121.840 337.830 122.055 ;
        RECT 338.000 121.885 338.690 122.055 ;
        RECT 335.780 121.525 336.635 121.605 ;
        RECT 331.360 120.825 331.630 121.315 ;
        RECT 331.800 120.115 331.970 121.315 ;
        RECT 332.640 120.825 332.910 121.315 ;
        RECT 333.240 121.145 333.690 121.315 ;
        RECT 333.240 120.825 333.410 121.145 ;
        RECT 332.140 120.285 333.650 120.635 ;
        RECT 334.080 120.115 334.250 121.315 ;
        RECT 334.520 120.825 334.790 121.315 ;
        RECT 334.960 120.115 335.130 121.315 ;
        RECT 335.865 120.115 336.035 121.315 ;
        RECT 336.305 120.825 336.475 121.315 ;
        RECT 336.745 120.115 336.915 121.315 ;
        RECT 337.560 120.115 337.730 121.315 ;
        RECT 338.000 120.825 338.170 121.885 ;
        RECT 340.000 121.840 340.330 122.055 ;
        RECT 340.500 121.885 341.190 122.055 ;
        RECT 338.340 121.485 338.670 121.655 ;
        RECT 338.440 120.115 338.610 121.315 ;
        RECT 339.180 120.115 339.570 121.480 ;
        RECT 340.060 120.115 340.230 121.315 ;
        RECT 340.500 120.825 340.670 121.885 ;
        RECT 340.840 121.485 341.170 121.655 ;
        RECT 340.940 120.115 341.110 121.315 ;
        RECT 341.780 120.435 341.950 122.250 ;
        RECT 342.240 122.225 342.630 123.165 ;
        RECT 343.080 122.225 343.250 123.875 ;
        RECT 343.580 123.380 343.910 123.550 ;
        RECT 343.640 122.225 343.910 123.165 ;
        RECT 344.080 122.225 344.250 123.875 ;
        RECT 342.120 121.605 342.290 121.935 ;
        RECT 342.460 121.855 342.630 122.225 ;
        RECT 343.740 121.935 343.910 122.225 ;
        RECT 344.520 121.935 344.690 123.165 ;
        RECT 345.080 122.225 345.250 123.875 ;
        RECT 345.520 122.225 345.790 123.165 ;
        RECT 345.960 122.225 346.130 123.875 ;
        RECT 342.460 121.685 343.570 121.855 ;
        RECT 342.460 121.315 342.630 121.685 ;
        RECT 343.740 121.610 344.350 121.935 ;
        RECT 343.740 121.315 343.910 121.610 ;
        RECT 344.180 121.605 344.350 121.610 ;
        RECT 344.520 121.605 345.450 121.935 ;
        RECT 344.520 121.315 344.690 121.605 ;
        RECT 345.620 121.315 345.790 122.225 ;
        RECT 342.360 120.825 342.630 121.315 ;
        RECT 342.800 120.115 342.970 121.315 ;
        RECT 343.640 120.825 343.910 121.315 ;
        RECT 344.240 121.145 344.690 121.315 ;
        RECT 344.240 120.825 344.410 121.145 ;
        RECT 343.140 120.285 344.650 120.635 ;
        RECT 345.080 120.115 345.250 121.315 ;
        RECT 345.520 120.825 345.790 121.315 ;
        RECT 345.960 120.115 346.130 121.315 ;
        RECT 298.500 119.865 346.500 120.115 ;
        RECT 298.500 117.625 346.000 117.875 ;
        RECT 298.865 115.975 299.035 117.625 ;
        RECT 299.305 115.975 299.475 116.915 ;
        RECT 299.745 115.975 299.915 117.625 ;
        RECT 300.430 116.035 300.820 117.625 ;
        RECT 301.280 116.500 301.450 117.330 ;
        RECT 301.820 117.130 302.150 117.300 ;
        RECT 301.280 116.000 301.570 116.500 ;
        RECT 298.780 115.685 299.635 115.765 ;
        RECT 298.750 115.355 299.635 115.685 ;
        RECT 298.780 115.275 299.635 115.355 ;
        RECT 298.865 113.865 299.035 115.065 ;
        RECT 299.305 114.575 299.475 115.065 ;
        RECT 299.745 113.865 299.915 115.065 ;
        RECT 300.430 113.865 300.820 115.230 ;
        RECT 301.280 114.185 301.450 116.000 ;
        RECT 301.740 115.975 302.130 116.915 ;
        RECT 302.580 115.975 302.750 117.625 ;
        RECT 303.080 117.130 303.410 117.300 ;
        RECT 303.140 115.975 303.410 116.915 ;
        RECT 303.580 115.975 303.750 117.625 ;
        RECT 301.620 115.355 301.790 115.685 ;
        RECT 301.960 115.605 302.130 115.975 ;
        RECT 303.240 115.685 303.410 115.975 ;
        RECT 304.020 115.685 304.190 116.915 ;
        RECT 304.580 115.975 304.750 117.625 ;
        RECT 305.020 115.975 305.290 116.915 ;
        RECT 305.460 115.975 305.630 117.625 ;
        RECT 306.180 116.035 306.570 117.625 ;
        RECT 306.930 116.035 307.320 117.625 ;
        RECT 307.680 116.035 308.070 117.625 ;
        RECT 308.280 116.500 308.450 117.330 ;
        RECT 308.820 117.130 309.150 117.300 ;
        RECT 308.280 116.000 308.570 116.500 ;
        RECT 301.960 115.435 303.070 115.605 ;
        RECT 301.960 115.065 302.130 115.435 ;
        RECT 303.240 115.360 303.850 115.685 ;
        RECT 303.240 115.065 303.410 115.360 ;
        RECT 303.680 115.355 303.850 115.360 ;
        RECT 304.020 115.355 304.950 115.685 ;
        RECT 304.020 115.065 304.190 115.355 ;
        RECT 305.120 115.065 305.290 115.975 ;
        RECT 301.860 114.575 302.130 115.065 ;
        RECT 302.300 113.865 302.470 115.065 ;
        RECT 303.140 114.575 303.410 115.065 ;
        RECT 303.740 114.895 304.190 115.065 ;
        RECT 303.740 114.575 303.910 114.895 ;
        RECT 302.640 114.035 304.150 114.385 ;
        RECT 304.580 113.865 304.750 115.065 ;
        RECT 305.020 114.575 305.290 115.065 ;
        RECT 305.460 113.865 305.630 115.065 ;
        RECT 306.180 113.865 306.570 115.230 ;
        RECT 306.930 113.865 307.320 115.230 ;
        RECT 307.680 113.865 308.070 115.230 ;
        RECT 308.280 114.185 308.450 116.000 ;
        RECT 308.740 115.975 309.130 116.915 ;
        RECT 309.580 115.975 309.750 117.625 ;
        RECT 310.080 117.130 310.410 117.300 ;
        RECT 310.140 115.975 310.410 116.915 ;
        RECT 310.580 115.975 310.750 117.625 ;
        RECT 308.620 115.355 308.790 115.685 ;
        RECT 308.960 115.605 309.130 115.975 ;
        RECT 310.240 115.685 310.410 115.975 ;
        RECT 311.020 115.685 311.190 116.915 ;
        RECT 311.580 115.975 311.750 117.625 ;
        RECT 312.020 115.975 312.290 116.915 ;
        RECT 312.460 115.975 312.630 117.625 ;
        RECT 313.180 116.035 313.570 117.625 ;
        RECT 313.930 116.035 314.320 117.625 ;
        RECT 314.865 115.975 315.035 117.625 ;
        RECT 315.305 115.975 315.475 116.915 ;
        RECT 315.745 115.975 315.915 117.625 ;
        RECT 316.430 116.035 316.820 117.625 ;
        RECT 317.280 116.500 317.450 117.330 ;
        RECT 317.820 117.130 318.150 117.300 ;
        RECT 317.280 116.000 317.570 116.500 ;
        RECT 308.960 115.435 310.070 115.605 ;
        RECT 308.960 115.065 309.130 115.435 ;
        RECT 310.240 115.360 310.850 115.685 ;
        RECT 310.240 115.065 310.410 115.360 ;
        RECT 310.680 115.355 310.850 115.360 ;
        RECT 311.020 115.355 311.950 115.685 ;
        RECT 311.020 115.065 311.190 115.355 ;
        RECT 312.120 115.065 312.290 115.975 ;
        RECT 314.780 115.685 315.635 115.765 ;
        RECT 314.750 115.355 315.635 115.685 ;
        RECT 314.780 115.275 315.635 115.355 ;
        RECT 308.860 114.575 309.130 115.065 ;
        RECT 309.300 113.865 309.470 115.065 ;
        RECT 310.140 114.575 310.410 115.065 ;
        RECT 310.740 114.895 311.190 115.065 ;
        RECT 310.740 114.575 310.910 114.895 ;
        RECT 309.640 114.035 311.150 114.385 ;
        RECT 311.580 113.865 311.750 115.065 ;
        RECT 312.020 114.575 312.290 115.065 ;
        RECT 312.460 113.865 312.630 115.065 ;
        RECT 313.180 113.865 313.570 115.230 ;
        RECT 313.930 113.865 314.320 115.230 ;
        RECT 314.865 113.865 315.035 115.065 ;
        RECT 315.305 114.575 315.475 115.065 ;
        RECT 315.745 113.865 315.915 115.065 ;
        RECT 316.430 113.865 316.820 115.230 ;
        RECT 317.280 114.185 317.450 116.000 ;
        RECT 317.740 115.975 318.130 116.915 ;
        RECT 318.580 115.975 318.750 117.625 ;
        RECT 319.080 117.130 319.410 117.300 ;
        RECT 319.140 115.975 319.410 116.915 ;
        RECT 319.580 115.975 319.750 117.625 ;
        RECT 317.620 115.355 317.790 115.685 ;
        RECT 317.960 115.605 318.130 115.975 ;
        RECT 319.240 115.685 319.410 115.975 ;
        RECT 320.020 115.685 320.190 116.915 ;
        RECT 320.580 115.975 320.750 117.625 ;
        RECT 321.020 115.975 321.290 116.915 ;
        RECT 321.460 115.975 321.630 117.625 ;
        RECT 322.030 116.500 322.200 117.330 ;
        RECT 322.570 117.130 322.900 117.300 ;
        RECT 322.030 116.000 322.320 116.500 ;
        RECT 317.960 115.435 319.070 115.605 ;
        RECT 317.960 115.065 318.130 115.435 ;
        RECT 319.240 115.360 319.850 115.685 ;
        RECT 319.240 115.065 319.410 115.360 ;
        RECT 319.680 115.355 319.850 115.360 ;
        RECT 320.020 115.355 320.950 115.685 ;
        RECT 320.020 115.065 320.190 115.355 ;
        RECT 321.120 115.065 321.290 115.975 ;
        RECT 317.860 114.575 318.130 115.065 ;
        RECT 318.300 113.865 318.470 115.065 ;
        RECT 319.140 114.575 319.410 115.065 ;
        RECT 319.740 114.895 320.190 115.065 ;
        RECT 319.740 114.575 319.910 114.895 ;
        RECT 318.640 114.035 320.150 114.385 ;
        RECT 320.580 113.865 320.750 115.065 ;
        RECT 321.020 114.575 321.290 115.065 ;
        RECT 321.460 113.865 321.630 115.065 ;
        RECT 322.030 114.185 322.200 116.000 ;
        RECT 322.490 115.975 322.880 116.915 ;
        RECT 323.330 115.975 323.500 117.625 ;
        RECT 323.830 117.130 324.160 117.300 ;
        RECT 323.890 115.975 324.160 116.915 ;
        RECT 324.330 115.975 324.500 117.625 ;
        RECT 322.370 115.355 322.540 115.685 ;
        RECT 322.710 115.605 322.880 115.975 ;
        RECT 323.990 115.685 324.160 115.975 ;
        RECT 324.770 115.685 324.940 116.915 ;
        RECT 325.330 115.975 325.500 117.625 ;
        RECT 325.770 115.975 326.040 116.915 ;
        RECT 326.210 115.975 326.380 117.625 ;
        RECT 326.930 116.035 327.320 117.625 ;
        RECT 327.865 115.975 328.035 117.625 ;
        RECT 328.305 115.975 328.475 116.915 ;
        RECT 328.745 115.975 328.915 117.625 ;
        RECT 329.365 115.975 329.535 117.625 ;
        RECT 329.805 115.975 329.975 116.915 ;
        RECT 330.245 115.975 330.415 117.625 ;
        RECT 330.865 115.975 331.035 117.625 ;
        RECT 331.305 115.975 331.475 116.915 ;
        RECT 331.745 115.975 331.915 117.625 ;
        RECT 332.430 116.035 332.820 117.625 ;
        RECT 333.280 116.500 333.450 117.330 ;
        RECT 333.820 117.130 334.150 117.300 ;
        RECT 333.280 116.000 333.570 116.500 ;
        RECT 322.710 115.435 323.820 115.605 ;
        RECT 322.710 115.065 322.880 115.435 ;
        RECT 323.990 115.360 324.600 115.685 ;
        RECT 323.990 115.065 324.160 115.360 ;
        RECT 324.430 115.355 324.600 115.360 ;
        RECT 324.770 115.355 325.700 115.685 ;
        RECT 324.770 115.065 324.940 115.355 ;
        RECT 325.870 115.065 326.040 115.975 ;
        RECT 327.780 115.685 328.635 115.765 ;
        RECT 329.280 115.685 330.135 115.765 ;
        RECT 330.780 115.685 331.635 115.765 ;
        RECT 327.750 115.355 328.635 115.685 ;
        RECT 329.250 115.355 330.135 115.685 ;
        RECT 330.750 115.355 331.635 115.685 ;
        RECT 327.780 115.275 328.635 115.355 ;
        RECT 329.280 115.275 330.135 115.355 ;
        RECT 330.780 115.275 331.635 115.355 ;
        RECT 322.610 114.575 322.880 115.065 ;
        RECT 323.050 113.865 323.220 115.065 ;
        RECT 323.890 114.575 324.160 115.065 ;
        RECT 324.490 114.895 324.940 115.065 ;
        RECT 324.490 114.575 324.660 114.895 ;
        RECT 323.390 114.035 324.900 114.385 ;
        RECT 325.330 113.865 325.500 115.065 ;
        RECT 325.770 114.575 326.040 115.065 ;
        RECT 326.210 113.865 326.380 115.065 ;
        RECT 326.930 113.865 327.320 115.230 ;
        RECT 327.865 113.865 328.035 115.065 ;
        RECT 328.305 114.575 328.475 115.065 ;
        RECT 328.745 113.865 328.915 115.065 ;
        RECT 329.365 113.865 329.535 115.065 ;
        RECT 329.805 114.575 329.975 115.065 ;
        RECT 330.245 113.865 330.415 115.065 ;
        RECT 330.865 113.865 331.035 115.065 ;
        RECT 331.305 114.575 331.475 115.065 ;
        RECT 331.745 113.865 331.915 115.065 ;
        RECT 332.430 113.865 332.820 115.230 ;
        RECT 333.280 114.185 333.450 116.000 ;
        RECT 333.740 115.975 334.130 116.915 ;
        RECT 334.580 115.975 334.750 117.625 ;
        RECT 335.080 117.130 335.410 117.300 ;
        RECT 335.140 115.975 335.410 116.915 ;
        RECT 335.580 115.975 335.750 117.625 ;
        RECT 333.620 115.355 333.790 115.685 ;
        RECT 333.960 115.605 334.130 115.975 ;
        RECT 335.240 115.685 335.410 115.975 ;
        RECT 336.020 115.685 336.190 116.915 ;
        RECT 336.580 115.975 336.750 117.625 ;
        RECT 337.020 115.975 337.290 116.915 ;
        RECT 337.460 115.975 337.630 117.625 ;
        RECT 338.180 116.035 338.570 117.625 ;
        RECT 338.930 116.035 339.320 117.625 ;
        RECT 339.780 116.500 339.950 117.330 ;
        RECT 340.320 117.130 340.650 117.300 ;
        RECT 339.780 116.000 340.070 116.500 ;
        RECT 333.960 115.435 335.070 115.605 ;
        RECT 333.960 115.065 334.130 115.435 ;
        RECT 335.240 115.360 335.850 115.685 ;
        RECT 335.240 115.065 335.410 115.360 ;
        RECT 335.680 115.355 335.850 115.360 ;
        RECT 336.020 115.355 336.950 115.685 ;
        RECT 336.020 115.065 336.190 115.355 ;
        RECT 337.120 115.065 337.290 115.975 ;
        RECT 333.860 114.575 334.130 115.065 ;
        RECT 334.300 113.865 334.470 115.065 ;
        RECT 335.140 114.575 335.410 115.065 ;
        RECT 335.740 114.895 336.190 115.065 ;
        RECT 335.740 114.575 335.910 114.895 ;
        RECT 334.640 114.035 336.150 114.385 ;
        RECT 336.580 113.865 336.750 115.065 ;
        RECT 337.020 114.575 337.290 115.065 ;
        RECT 337.460 113.865 337.630 115.065 ;
        RECT 338.180 113.865 338.570 115.230 ;
        RECT 338.930 113.865 339.320 115.230 ;
        RECT 339.780 114.185 339.950 116.000 ;
        RECT 340.240 115.975 340.630 116.915 ;
        RECT 341.080 115.975 341.250 117.625 ;
        RECT 341.580 117.130 341.910 117.300 ;
        RECT 341.640 115.975 341.910 116.915 ;
        RECT 342.080 115.975 342.250 117.625 ;
        RECT 340.120 115.355 340.290 115.685 ;
        RECT 340.460 115.605 340.630 115.975 ;
        RECT 341.740 115.685 341.910 115.975 ;
        RECT 342.520 115.685 342.690 116.915 ;
        RECT 343.080 115.975 343.250 117.625 ;
        RECT 343.520 115.975 343.790 116.915 ;
        RECT 343.960 115.975 344.130 117.625 ;
        RECT 344.680 116.035 345.070 117.625 ;
        RECT 345.430 116.035 345.820 117.625 ;
        RECT 340.460 115.435 341.570 115.605 ;
        RECT 340.460 115.065 340.630 115.435 ;
        RECT 341.740 115.360 342.350 115.685 ;
        RECT 341.740 115.065 341.910 115.360 ;
        RECT 342.180 115.355 342.350 115.360 ;
        RECT 342.520 115.355 343.450 115.685 ;
        RECT 342.520 115.065 342.690 115.355 ;
        RECT 343.620 115.065 343.790 115.975 ;
        RECT 340.360 114.575 340.630 115.065 ;
        RECT 340.800 113.865 340.970 115.065 ;
        RECT 341.640 114.575 341.910 115.065 ;
        RECT 342.240 114.895 342.690 115.065 ;
        RECT 342.240 114.575 342.410 114.895 ;
        RECT 341.140 114.035 342.650 114.385 ;
        RECT 343.080 113.865 343.250 115.065 ;
        RECT 343.520 114.575 343.790 115.065 ;
        RECT 343.960 113.865 344.130 115.065 ;
        RECT 344.680 113.865 345.070 115.230 ;
        RECT 345.430 113.865 345.820 115.230 ;
        RECT 298.500 113.615 346.000 113.865 ;
        RECT 349.750 112.750 350.250 125.750 ;
        RECT 388.125 123.875 388.375 127.375 ;
        RECT 389.665 126.500 389.835 127.000 ;
        RECT 388.780 125.230 389.260 126.270 ;
        RECT 389.530 125.230 389.970 126.270 ;
        RECT 390.240 125.230 390.720 126.270 ;
        RECT 389.665 124.500 389.835 125.000 ;
        RECT 391.125 123.875 391.375 127.375 ;
        RECT 388.125 123.625 391.375 123.875 ;
        RECT 388.125 120.125 388.375 123.625 ;
        RECT 389.665 122.750 389.835 123.250 ;
        RECT 388.780 121.480 389.260 122.520 ;
        RECT 389.530 121.480 389.970 122.520 ;
        RECT 390.240 121.480 390.720 122.520 ;
        RECT 389.665 120.750 389.835 121.250 ;
        RECT 391.125 120.125 391.375 123.625 ;
        RECT 388.125 119.875 391.375 120.125 ;
        RECT 397.625 149.875 400.875 150.125 ;
        RECT 397.625 146.375 397.875 149.875 ;
        RECT 399.165 149.000 399.335 149.500 ;
        RECT 398.280 147.730 398.760 148.770 ;
        RECT 399.030 147.730 399.470 148.770 ;
        RECT 399.740 147.730 400.220 148.770 ;
        RECT 399.165 147.000 399.335 147.500 ;
        RECT 400.625 146.375 400.875 149.875 ;
        RECT 397.625 146.125 400.875 146.375 ;
        RECT 397.625 142.625 397.875 146.125 ;
        RECT 399.165 145.250 399.335 145.750 ;
        RECT 398.280 143.980 398.760 145.020 ;
        RECT 399.030 143.980 399.470 145.020 ;
        RECT 399.740 143.980 400.220 145.020 ;
        RECT 399.165 143.250 399.335 143.750 ;
        RECT 400.625 142.625 400.875 146.125 ;
        RECT 397.625 142.375 400.875 142.625 ;
        RECT 397.625 138.875 397.875 142.375 ;
        RECT 399.165 141.500 399.335 142.000 ;
        RECT 398.280 140.230 398.760 141.270 ;
        RECT 399.030 140.230 399.470 141.270 ;
        RECT 399.740 140.230 400.220 141.270 ;
        RECT 399.165 139.500 399.335 140.000 ;
        RECT 400.625 138.875 400.875 142.375 ;
        RECT 397.625 138.625 400.875 138.875 ;
        RECT 397.625 135.125 397.875 138.625 ;
        RECT 399.165 137.750 399.335 138.250 ;
        RECT 398.280 136.480 398.760 137.520 ;
        RECT 399.030 136.480 399.470 137.520 ;
        RECT 399.740 136.480 400.220 137.520 ;
        RECT 399.165 135.750 399.335 136.250 ;
        RECT 400.625 135.125 400.875 138.625 ;
        RECT 397.625 134.875 400.875 135.125 ;
        RECT 397.625 131.375 397.875 134.875 ;
        RECT 399.165 134.000 399.335 134.500 ;
        RECT 398.280 132.730 398.760 133.770 ;
        RECT 399.030 132.730 399.470 133.770 ;
        RECT 399.740 132.730 400.220 133.770 ;
        RECT 399.165 132.000 399.335 132.500 ;
        RECT 400.625 131.375 400.875 134.875 ;
        RECT 397.625 131.125 400.875 131.375 ;
        RECT 397.625 127.625 397.875 131.125 ;
        RECT 399.165 130.250 399.335 130.750 ;
        RECT 398.280 128.980 398.760 130.020 ;
        RECT 399.030 128.980 399.470 130.020 ;
        RECT 399.740 128.980 400.220 130.020 ;
        RECT 399.165 128.250 399.335 128.750 ;
        RECT 400.625 127.625 400.875 131.125 ;
        RECT 397.625 127.375 400.875 127.625 ;
        RECT 397.625 123.875 397.875 127.375 ;
        RECT 399.165 126.500 399.335 127.000 ;
        RECT 398.280 125.230 398.760 126.270 ;
        RECT 399.030 125.230 399.470 126.270 ;
        RECT 399.740 125.230 400.220 126.270 ;
        RECT 399.165 124.500 399.335 125.000 ;
        RECT 400.625 123.875 400.875 127.375 ;
        RECT 397.625 123.625 400.875 123.875 ;
        RECT 397.625 120.125 397.875 123.625 ;
        RECT 399.165 122.750 399.335 123.250 ;
        RECT 398.280 121.480 398.760 122.520 ;
        RECT 399.030 121.480 399.470 122.520 ;
        RECT 399.740 121.480 400.220 122.520 ;
        RECT 399.165 120.750 399.335 121.250 ;
        RECT 400.625 120.125 400.875 123.625 ;
        RECT 397.625 119.875 400.875 120.125 ;
        RECT 407.125 149.875 410.375 150.125 ;
        RECT 407.125 146.375 407.375 149.875 ;
        RECT 408.665 149.000 408.835 149.500 ;
        RECT 407.780 147.730 408.260 148.770 ;
        RECT 408.530 147.730 408.970 148.770 ;
        RECT 409.240 147.730 409.720 148.770 ;
        RECT 408.665 147.000 408.835 147.500 ;
        RECT 410.125 146.375 410.375 149.875 ;
        RECT 407.125 146.125 410.375 146.375 ;
        RECT 407.125 142.625 407.375 146.125 ;
        RECT 408.665 145.250 408.835 145.750 ;
        RECT 407.780 143.980 408.260 145.020 ;
        RECT 408.530 143.980 408.970 145.020 ;
        RECT 409.240 143.980 409.720 145.020 ;
        RECT 408.665 143.250 408.835 143.750 ;
        RECT 410.125 142.625 410.375 146.125 ;
        RECT 407.125 142.375 410.375 142.625 ;
        RECT 407.125 138.875 407.375 142.375 ;
        RECT 408.665 141.500 408.835 142.000 ;
        RECT 407.780 140.230 408.260 141.270 ;
        RECT 408.530 140.230 408.970 141.270 ;
        RECT 409.240 140.230 409.720 141.270 ;
        RECT 408.665 139.500 408.835 140.000 ;
        RECT 410.125 138.875 410.375 142.375 ;
        RECT 407.125 138.625 410.375 138.875 ;
        RECT 407.125 135.125 407.375 138.625 ;
        RECT 408.665 137.750 408.835 138.250 ;
        RECT 407.780 136.480 408.260 137.520 ;
        RECT 408.530 136.480 408.970 137.520 ;
        RECT 409.240 136.480 409.720 137.520 ;
        RECT 408.665 135.750 408.835 136.250 ;
        RECT 410.125 135.125 410.375 138.625 ;
        RECT 407.125 134.875 410.375 135.125 ;
        RECT 407.125 131.375 407.375 134.875 ;
        RECT 408.665 134.000 408.835 134.500 ;
        RECT 407.780 132.730 408.260 133.770 ;
        RECT 408.530 132.730 408.970 133.770 ;
        RECT 409.240 132.730 409.720 133.770 ;
        RECT 408.665 132.000 408.835 132.500 ;
        RECT 410.125 131.375 410.375 134.875 ;
        RECT 407.125 131.125 410.375 131.375 ;
        RECT 407.125 127.625 407.375 131.125 ;
        RECT 408.665 130.250 408.835 130.750 ;
        RECT 407.780 128.980 408.260 130.020 ;
        RECT 408.530 128.980 408.970 130.020 ;
        RECT 409.240 128.980 409.720 130.020 ;
        RECT 408.665 128.250 408.835 128.750 ;
        RECT 410.125 127.625 410.375 131.125 ;
        RECT 407.125 127.375 410.375 127.625 ;
        RECT 407.125 123.875 407.375 127.375 ;
        RECT 408.665 126.500 408.835 127.000 ;
        RECT 407.780 125.230 408.260 126.270 ;
        RECT 408.530 125.230 408.970 126.270 ;
        RECT 409.240 125.230 409.720 126.270 ;
        RECT 408.665 124.500 408.835 125.000 ;
        RECT 410.125 123.875 410.375 127.375 ;
        RECT 407.125 123.625 410.375 123.875 ;
        RECT 407.125 120.125 407.375 123.625 ;
        RECT 408.665 122.750 408.835 123.250 ;
        RECT 407.780 121.480 408.260 122.520 ;
        RECT 408.530 121.480 408.970 122.520 ;
        RECT 409.240 121.480 409.720 122.520 ;
        RECT 408.665 120.750 408.835 121.250 ;
        RECT 410.125 120.125 410.375 123.625 ;
        RECT 407.125 119.875 410.375 120.125 ;
        RECT 294.250 112.250 350.250 112.750 ;
      LAYER met1 ;
        RECT 288.500 205.000 427.000 209.000 ;
        RECT 288.500 200.000 425.000 204.000 ;
        RECT 322.750 197.750 348.250 199.000 ;
        RECT 325.750 193.000 326.250 197.750 ;
        RECT 326.525 197.000 328.520 197.500 ;
        RECT 328.935 197.000 330.925 197.750 ;
        RECT 326.525 194.640 326.755 197.000 ;
        RECT 326.965 194.500 327.195 196.640 ;
        RECT 327.405 194.640 327.635 197.000 ;
        RECT 327.845 194.500 328.075 196.640 ;
        RECT 328.285 194.640 328.515 197.000 ;
        RECT 328.935 194.640 329.165 197.000 ;
        RECT 326.520 194.000 328.075 194.500 ;
        RECT 329.375 194.500 329.605 196.640 ;
        RECT 329.815 194.640 330.045 197.000 ;
        RECT 330.255 194.500 330.485 196.640 ;
        RECT 330.695 194.640 330.925 197.000 ;
        RECT 331.345 197.000 333.335 197.750 ;
        RECT 331.345 194.640 331.575 197.000 ;
        RECT 331.785 194.500 332.015 196.640 ;
        RECT 332.225 194.640 332.455 197.000 ;
        RECT 332.665 194.500 332.895 196.640 ;
        RECT 333.105 194.640 333.335 197.000 ;
        RECT 333.755 197.000 335.745 197.750 ;
        RECT 333.755 194.640 333.985 197.000 ;
        RECT 334.195 194.500 334.425 196.640 ;
        RECT 334.635 194.640 334.865 197.000 ;
        RECT 335.075 194.500 335.305 196.640 ;
        RECT 335.515 194.640 335.745 197.000 ;
        RECT 336.165 197.000 338.160 197.500 ;
        RECT 338.575 197.000 340.565 197.750 ;
        RECT 336.165 194.640 336.395 197.000 ;
        RECT 336.605 194.500 336.835 196.640 ;
        RECT 337.045 194.640 337.275 197.000 ;
        RECT 337.485 194.500 337.715 196.640 ;
        RECT 337.925 194.640 338.155 197.000 ;
        RECT 338.575 194.640 338.805 197.000 ;
        RECT 339.015 194.500 339.245 196.640 ;
        RECT 339.455 194.640 339.685 197.000 ;
        RECT 339.895 194.500 340.125 196.640 ;
        RECT 340.335 194.640 340.565 197.000 ;
        RECT 340.985 197.000 342.975 197.750 ;
        RECT 340.985 194.640 341.215 197.000 ;
        RECT 341.425 194.500 341.655 196.640 ;
        RECT 341.865 194.640 342.095 197.000 ;
        RECT 342.305 194.500 342.535 196.640 ;
        RECT 342.745 194.640 342.975 197.000 ;
        RECT 329.375 194.000 330.930 194.500 ;
        RECT 331.340 194.000 332.895 194.500 ;
        RECT 333.750 194.000 335.750 194.500 ;
        RECT 336.160 194.000 337.715 194.500 ;
        RECT 338.570 194.000 340.125 194.500 ;
        RECT 340.980 194.000 342.535 194.500 ;
        RECT 327.270 193.250 330.180 193.750 ;
        RECT 330.430 193.250 332.590 193.750 ;
        RECT 334.500 193.250 335.000 193.750 ;
        RECT 336.910 193.250 339.070 193.750 ;
        RECT 339.320 193.250 342.230 193.750 ;
        RECT 343.250 193.000 343.750 197.750 ;
        RECT 382.750 196.000 411.250 197.000 ;
        RECT 322.750 192.500 348.250 193.000 ;
        RECT 349.250 192.750 355.750 194.000 ;
        RECT 387.500 193.000 388.500 196.000 ;
        RECT 388.750 195.000 389.250 195.500 ;
        RECT 389.500 195.250 390.000 195.750 ;
        RECT 390.250 195.000 390.750 195.500 ;
        RECT 388.750 194.000 389.290 195.000 ;
        RECT 389.500 194.000 390.000 195.000 ;
        RECT 390.210 194.000 390.750 195.000 ;
        RECT 389.500 193.250 390.000 193.750 ;
        RECT 391.000 193.000 392.000 196.000 ;
        RECT 324.250 191.750 327.770 192.250 ;
        RECT 328.020 191.750 341.480 192.250 ;
        RECT 341.730 191.750 345.250 192.250 ;
        RECT 326.520 191.000 336.660 191.500 ;
        RECT 324.250 190.250 327.770 190.750 ;
        RECT 331.340 190.250 341.480 190.750 ;
        RECT 341.730 190.250 345.250 190.750 ;
        RECT 328.020 189.500 338.160 190.000 ;
        RECT 349.250 189.750 349.750 192.750 ;
        RECT 350.750 192.000 351.250 192.500 ;
        RECT 350.000 190.750 350.895 191.750 ;
        RECT 351.105 190.750 352.000 191.750 ;
        RECT 350.750 190.000 351.250 190.500 ;
        RECT 352.250 189.750 352.750 192.750 ;
        RECT 353.750 192.000 354.250 192.500 ;
        RECT 353.000 190.750 353.895 191.750 ;
        RECT 354.105 190.750 355.000 191.750 ;
        RECT 353.750 190.000 354.250 190.500 ;
        RECT 355.250 189.750 355.750 192.750 ;
        RECT 374.500 192.500 381.750 193.000 ;
        RECT 387.500 192.500 392.000 193.000 ;
        RECT 349.250 189.250 355.750 189.750 ;
        RECT 387.500 189.250 388.500 192.500 ;
        RECT 388.750 191.250 389.250 191.750 ;
        RECT 389.500 191.500 390.000 192.000 ;
        RECT 390.250 191.250 390.750 191.750 ;
        RECT 388.750 190.250 389.290 191.250 ;
        RECT 389.500 190.250 390.000 191.250 ;
        RECT 390.210 190.250 390.750 191.250 ;
        RECT 389.500 189.500 390.000 190.000 ;
        RECT 391.000 189.250 392.000 192.500 ;
        RECT 321.250 188.750 346.750 189.250 ;
        RECT 372.500 188.750 381.750 189.250 ;
        RECT 387.500 188.750 392.000 189.250 ;
        RECT 325.750 184.750 326.250 188.750 ;
        RECT 327.270 188.000 330.180 188.500 ;
        RECT 330.430 188.000 332.590 188.500 ;
        RECT 334.500 188.000 335.000 188.500 ;
        RECT 336.910 188.000 339.070 188.500 ;
        RECT 339.320 188.000 342.230 188.500 ;
        RECT 326.520 187.250 328.075 187.750 ;
        RECT 326.525 185.500 326.755 187.110 ;
        RECT 326.965 186.110 327.195 187.250 ;
        RECT 327.405 185.500 327.635 187.110 ;
        RECT 327.845 186.110 328.075 187.250 ;
        RECT 329.375 187.250 330.930 187.750 ;
        RECT 331.785 187.250 333.340 187.750 ;
        RECT 333.750 187.250 335.750 187.750 ;
        RECT 336.605 187.250 338.160 187.750 ;
        RECT 338.570 187.250 340.125 187.750 ;
        RECT 340.980 187.250 342.535 187.750 ;
        RECT 328.285 185.500 328.515 187.110 ;
        RECT 328.935 185.500 329.165 187.110 ;
        RECT 329.375 186.110 329.605 187.250 ;
        RECT 329.815 185.500 330.045 187.110 ;
        RECT 330.255 186.110 330.485 187.250 ;
        RECT 330.695 185.500 330.925 187.110 ;
        RECT 331.345 185.500 331.575 187.110 ;
        RECT 331.785 186.110 332.015 187.250 ;
        RECT 332.225 185.500 332.455 187.110 ;
        RECT 332.665 186.110 332.895 187.250 ;
        RECT 333.105 185.500 333.335 187.110 ;
        RECT 326.525 185.000 328.520 185.500 ;
        RECT 328.935 184.750 330.925 185.500 ;
        RECT 331.340 185.000 333.335 185.500 ;
        RECT 333.755 185.500 333.985 187.110 ;
        RECT 334.195 186.110 334.425 187.250 ;
        RECT 334.635 185.500 334.865 187.110 ;
        RECT 335.075 186.110 335.305 187.250 ;
        RECT 335.515 185.500 335.745 187.110 ;
        RECT 333.755 184.750 335.745 185.500 ;
        RECT 336.165 185.500 336.395 187.110 ;
        RECT 336.605 186.110 336.835 187.250 ;
        RECT 337.045 185.500 337.275 187.110 ;
        RECT 337.485 186.110 337.715 187.250 ;
        RECT 337.925 185.500 338.155 187.110 ;
        RECT 336.165 184.750 338.155 185.500 ;
        RECT 338.575 185.500 338.805 187.110 ;
        RECT 339.015 186.110 339.245 187.250 ;
        RECT 339.455 185.500 339.685 187.110 ;
        RECT 339.895 186.110 340.125 187.250 ;
        RECT 340.335 185.500 340.565 187.110 ;
        RECT 338.575 184.750 340.565 185.500 ;
        RECT 340.985 185.500 341.215 187.110 ;
        RECT 341.425 186.110 341.655 187.250 ;
        RECT 341.865 185.500 342.095 187.110 ;
        RECT 342.305 186.110 342.535 187.250 ;
        RECT 342.745 185.500 342.975 187.110 ;
        RECT 340.985 184.750 342.975 185.500 ;
        RECT 343.250 184.750 343.750 188.750 ;
        RECT 387.500 185.500 388.500 188.750 ;
        RECT 388.750 187.500 389.250 188.000 ;
        RECT 389.500 187.750 390.000 188.250 ;
        RECT 390.250 187.500 390.750 188.000 ;
        RECT 388.750 186.500 389.290 187.500 ;
        RECT 389.500 186.500 390.000 187.500 ;
        RECT 390.210 186.500 390.750 187.500 ;
        RECT 389.500 185.750 390.000 186.250 ;
        RECT 391.000 185.500 392.000 188.750 ;
        RECT 370.500 185.000 381.750 185.500 ;
        RECT 387.500 185.000 392.000 185.500 ;
        RECT 290.000 183.120 320.500 183.600 ;
        RECT 321.250 183.500 346.750 184.750 ;
        RECT 387.500 181.750 388.500 185.000 ;
        RECT 388.750 183.750 389.250 184.250 ;
        RECT 389.500 184.000 390.000 184.500 ;
        RECT 390.250 183.750 390.750 184.250 ;
        RECT 388.750 182.750 389.290 183.750 ;
        RECT 389.500 182.750 390.000 183.750 ;
        RECT 390.210 182.750 390.750 183.750 ;
        RECT 389.500 182.000 390.000 182.500 ;
        RECT 391.000 181.750 392.000 185.000 ;
        RECT 368.500 181.250 381.750 181.750 ;
        RECT 387.500 181.250 392.000 181.750 ;
        RECT 291.500 180.400 320.500 180.880 ;
        RECT 312.410 180.000 312.730 180.260 ;
        RECT 312.870 180.000 313.190 180.260 ;
        RECT 310.570 179.860 310.890 179.920 ;
        RECT 313.345 179.860 313.635 179.905 ;
        RECT 310.570 179.720 313.635 179.860 ;
        RECT 310.570 179.660 310.890 179.720 ;
        RECT 313.345 179.675 313.635 179.720 ;
        RECT 297.230 179.520 297.550 179.580 ;
        RECT 299.070 179.520 299.390 179.580 ;
        RECT 311.030 179.520 311.350 179.580 ;
        RECT 311.505 179.520 311.795 179.565 ;
        RECT 297.230 179.380 311.795 179.520 ;
        RECT 297.230 179.320 297.550 179.380 ;
        RECT 299.070 179.320 299.390 179.380 ;
        RECT 311.030 179.320 311.350 179.380 ;
        RECT 311.505 179.335 311.795 179.380 ;
        RECT 299.990 178.980 300.310 179.240 ;
        RECT 314.250 178.840 314.570 178.900 ;
        RECT 314.710 178.840 315.030 178.900 ;
        RECT 314.250 178.700 315.030 178.840 ;
        RECT 314.250 178.640 314.570 178.700 ;
        RECT 314.710 178.640 315.030 178.700 ;
        RECT 298.150 178.300 298.470 178.560 ;
        RECT 290.000 177.680 320.500 178.160 ;
        RECT 387.500 178.000 388.500 181.250 ;
        RECT 388.750 180.000 389.250 180.500 ;
        RECT 389.500 180.250 390.000 180.750 ;
        RECT 390.250 180.000 390.750 180.500 ;
        RECT 388.750 179.000 389.290 180.000 ;
        RECT 389.500 179.000 390.000 180.000 ;
        RECT 390.210 179.000 390.750 180.000 ;
        RECT 389.500 178.250 390.000 178.750 ;
        RECT 391.000 178.000 392.000 181.250 ;
        RECT 300.465 177.280 300.785 177.540 ;
        RECT 312.870 177.480 313.190 177.540 ;
        RECT 366.500 177.500 381.750 178.000 ;
        RECT 387.500 177.500 392.000 178.000 ;
        RECT 310.660 177.340 313.190 177.480 ;
        RECT 299.990 177.140 300.310 177.200 ;
        RECT 310.660 177.140 310.800 177.340 ;
        RECT 299.990 177.000 310.800 177.140 ;
        RECT 299.990 176.940 300.310 177.000 ;
        RECT 311.030 176.940 311.350 177.200 ;
        RECT 311.580 177.185 311.720 177.340 ;
        RECT 312.870 177.280 313.190 177.340 ;
        RECT 311.505 176.955 311.795 177.185 ;
        RECT 296.770 176.800 297.090 176.860 ;
        RECT 311.120 176.800 311.260 176.940 ;
        RECT 312.425 176.800 312.715 176.845 ;
        RECT 296.770 176.660 300.220 176.800 ;
        RECT 311.120 176.660 312.715 176.800 ;
        RECT 296.770 176.600 297.090 176.660 ;
        RECT 296.310 176.460 296.630 176.520 ;
        RECT 297.690 176.460 298.010 176.520 ;
        RECT 300.080 176.505 300.220 176.660 ;
        RECT 312.425 176.615 312.715 176.660 ;
        RECT 299.085 176.460 299.375 176.505 ;
        RECT 296.310 176.320 297.460 176.460 ;
        RECT 296.310 176.260 296.630 176.320 ;
        RECT 295.850 175.920 296.170 176.180 ;
        RECT 296.770 175.920 297.090 176.180 ;
        RECT 297.320 176.120 297.460 176.320 ;
        RECT 297.690 176.320 299.375 176.460 ;
        RECT 297.690 176.260 298.010 176.320 ;
        RECT 299.085 176.275 299.375 176.320 ;
        RECT 300.005 176.275 300.295 176.505 ;
        RECT 311.045 176.275 311.335 176.505 ;
        RECT 298.150 176.120 298.470 176.180 ;
        RECT 298.625 176.120 298.915 176.165 ;
        RECT 297.320 175.980 297.920 176.120 ;
        RECT 297.230 175.580 297.550 175.840 ;
        RECT 297.780 175.825 297.920 175.980 ;
        RECT 298.150 175.980 298.915 176.120 ;
        RECT 298.150 175.920 298.470 175.980 ;
        RECT 298.625 175.935 298.915 175.980 ;
        RECT 311.120 176.120 311.260 176.275 ;
        RECT 312.410 176.120 312.730 176.180 ;
        RECT 311.120 175.980 312.730 176.120 ;
        RECT 297.705 175.780 297.995 175.825 ;
        RECT 311.120 175.780 311.260 175.980 ;
        RECT 312.410 175.920 312.730 175.980 ;
        RECT 297.705 175.640 311.260 175.780 ;
        RECT 312.870 175.780 313.190 175.840 ;
        RECT 313.330 175.780 313.650 175.840 ;
        RECT 312.870 175.640 313.650 175.780 ;
        RECT 297.705 175.595 297.995 175.640 ;
        RECT 312.870 175.580 313.190 175.640 ;
        RECT 313.330 175.580 313.650 175.640 ;
        RECT 291.500 174.960 320.500 175.440 ;
        RECT 296.270 174.620 297.230 174.760 ;
        RECT 387.500 174.250 388.500 177.500 ;
        RECT 388.750 176.250 389.250 176.750 ;
        RECT 389.500 176.500 390.000 177.000 ;
        RECT 390.250 176.250 390.750 176.750 ;
        RECT 388.750 175.250 389.290 176.250 ;
        RECT 389.500 175.250 390.000 176.250 ;
        RECT 390.210 175.250 390.750 176.250 ;
        RECT 389.500 174.500 390.000 175.000 ;
        RECT 391.000 174.250 392.000 177.500 ;
        RECT 295.865 174.080 296.155 174.125 ;
        RECT 297.230 174.080 297.550 174.140 ;
        RECT 299.530 174.080 299.850 174.140 ;
        RECT 295.865 173.940 299.850 174.080 ;
        RECT 295.865 173.895 296.155 173.940 ;
        RECT 297.230 173.880 297.550 173.940 ;
        RECT 299.530 173.880 299.850 173.940 ;
        RECT 296.310 173.540 296.630 173.800 ;
        RECT 364.500 173.750 381.750 174.250 ;
        RECT 387.500 173.750 392.000 174.250 ;
        RECT 298.610 173.400 298.930 173.460 ;
        RECT 299.990 173.400 300.310 173.460 ;
        RECT 296.860 173.260 300.310 173.400 ;
        RECT 296.860 173.105 297.000 173.260 ;
        RECT 298.610 173.200 298.930 173.260 ;
        RECT 299.990 173.200 300.310 173.260 ;
        RECT 296.785 172.875 297.075 173.105 ;
        RECT 297.690 172.860 298.010 173.120 ;
        RECT 290.000 172.240 320.500 172.720 ;
        RECT 296.770 171.700 297.090 171.760 ;
        RECT 299.085 171.700 299.375 171.745 ;
        RECT 296.770 171.560 299.375 171.700 ;
        RECT 296.770 171.500 297.090 171.560 ;
        RECT 299.085 171.515 299.375 171.560 ;
        RECT 297.690 171.360 298.010 171.420 ;
        RECT 298.150 171.360 298.470 171.420 ;
        RECT 297.690 171.220 298.470 171.360 ;
        RECT 297.690 171.160 298.010 171.220 ;
        RECT 298.150 171.160 298.470 171.220 ;
        RECT 299.545 170.835 299.835 171.065 ;
        RECT 311.030 171.020 311.350 171.080 ;
        RECT 311.965 171.020 312.255 171.065 ;
        RECT 311.030 170.880 312.255 171.020 ;
        RECT 296.310 170.680 296.630 170.740 ;
        RECT 298.150 170.680 298.470 170.740 ;
        RECT 299.620 170.680 299.760 170.835 ;
        RECT 311.030 170.820 311.350 170.880 ;
        RECT 311.965 170.835 312.255 170.880 ;
        RECT 312.870 170.820 313.190 171.080 ;
        RECT 296.310 170.540 299.760 170.680 ;
        RECT 310.570 170.680 310.890 170.740 ;
        RECT 311.505 170.680 311.795 170.725 ;
        RECT 310.570 170.540 311.795 170.680 ;
        RECT 296.310 170.480 296.630 170.540 ;
        RECT 298.150 170.480 298.470 170.540 ;
        RECT 310.570 170.480 310.890 170.540 ;
        RECT 311.505 170.495 311.795 170.540 ;
        RECT 313.805 170.680 314.095 170.725 ;
        RECT 317.010 170.680 317.330 170.740 ;
        RECT 313.805 170.540 317.330 170.680 ;
        RECT 313.805 170.495 314.095 170.540 ;
        RECT 317.010 170.480 317.330 170.540 ;
        RECT 387.500 170.500 388.500 173.750 ;
        RECT 388.750 172.500 389.250 173.000 ;
        RECT 389.500 172.750 390.000 173.250 ;
        RECT 390.250 172.500 390.750 173.000 ;
        RECT 388.750 171.500 389.290 172.500 ;
        RECT 389.500 171.500 390.000 172.500 ;
        RECT 390.210 171.500 390.750 172.500 ;
        RECT 389.500 170.750 390.000 171.250 ;
        RECT 391.000 170.500 392.000 173.750 ;
        RECT 295.390 170.340 295.710 170.400 ;
        RECT 297.245 170.340 297.535 170.385 ;
        RECT 295.390 170.200 297.535 170.340 ;
        RECT 295.390 170.140 295.710 170.200 ;
        RECT 297.245 170.155 297.535 170.200 ;
        RECT 362.500 170.000 381.750 170.500 ;
        RECT 387.500 170.000 392.000 170.500 ;
        RECT 291.500 169.520 320.500 170.000 ;
        RECT 311.030 168.640 311.350 168.700 ;
        RECT 312.425 168.640 312.715 168.685 ;
        RECT 311.030 168.500 312.715 168.640 ;
        RECT 311.030 168.440 311.350 168.500 ;
        RECT 312.425 168.455 312.715 168.500 ;
        RECT 313.330 167.760 313.650 168.020 ;
        RECT 290.000 166.800 320.500 167.280 ;
        RECT 387.500 166.750 388.500 170.000 ;
        RECT 388.750 168.750 389.250 169.250 ;
        RECT 389.500 169.000 390.000 169.500 ;
        RECT 390.250 168.750 390.750 169.250 ;
        RECT 388.750 167.750 389.290 168.750 ;
        RECT 389.500 167.750 390.000 168.750 ;
        RECT 390.210 167.750 390.750 168.750 ;
        RECT 389.500 167.000 390.000 167.500 ;
        RECT 391.000 166.750 392.000 170.000 ;
        RECT 298.610 166.600 298.930 166.660 ;
        RECT 301.845 166.600 302.135 166.645 ;
        RECT 298.610 166.460 302.135 166.600 ;
        RECT 298.610 166.400 298.930 166.460 ;
        RECT 301.845 166.415 302.135 166.460 ;
        RECT 312.885 166.600 313.175 166.645 ;
        RECT 314.250 166.600 314.570 166.660 ;
        RECT 312.885 166.460 314.570 166.600 ;
        RECT 312.885 166.415 313.175 166.460 ;
        RECT 297.230 165.920 297.550 165.980 ;
        RECT 297.705 165.920 297.995 165.965 ;
        RECT 301.415 165.920 301.735 165.980 ;
        RECT 297.230 165.780 301.735 165.920 ;
        RECT 301.920 165.920 302.060 166.415 ;
        RECT 314.250 166.400 314.570 166.460 ;
        RECT 360.500 166.250 381.750 166.750 ;
        RECT 387.500 166.250 392.000 166.750 ;
        RECT 397.000 193.000 398.000 196.000 ;
        RECT 398.250 195.000 398.750 195.500 ;
        RECT 399.000 195.250 399.500 195.750 ;
        RECT 399.750 195.000 400.250 195.500 ;
        RECT 398.250 194.000 398.790 195.000 ;
        RECT 399.000 194.000 399.500 195.000 ;
        RECT 399.710 194.000 400.250 195.000 ;
        RECT 399.000 193.250 399.500 193.750 ;
        RECT 400.500 193.000 401.500 196.000 ;
        RECT 397.000 192.500 401.500 193.000 ;
        RECT 397.000 189.250 398.000 192.500 ;
        RECT 398.250 191.250 398.750 191.750 ;
        RECT 399.000 191.500 399.500 192.000 ;
        RECT 399.750 191.250 400.250 191.750 ;
        RECT 398.250 190.250 398.790 191.250 ;
        RECT 399.000 190.250 399.500 191.250 ;
        RECT 399.710 190.250 400.250 191.250 ;
        RECT 399.000 189.500 399.500 190.000 ;
        RECT 400.500 189.250 401.500 192.500 ;
        RECT 397.000 188.750 401.500 189.250 ;
        RECT 397.000 185.500 398.000 188.750 ;
        RECT 398.250 187.500 398.750 188.000 ;
        RECT 399.000 187.750 399.500 188.250 ;
        RECT 399.750 187.500 400.250 188.000 ;
        RECT 398.250 186.500 398.790 187.500 ;
        RECT 399.000 186.500 399.500 187.500 ;
        RECT 399.710 186.500 400.250 187.500 ;
        RECT 399.000 185.750 399.500 186.250 ;
        RECT 400.500 185.500 401.500 188.750 ;
        RECT 397.000 185.000 401.500 185.500 ;
        RECT 397.000 181.750 398.000 185.000 ;
        RECT 398.250 183.750 398.750 184.250 ;
        RECT 399.000 184.000 399.500 184.500 ;
        RECT 399.750 183.750 400.250 184.250 ;
        RECT 398.250 182.750 398.790 183.750 ;
        RECT 399.000 182.750 399.500 183.750 ;
        RECT 399.710 182.750 400.250 183.750 ;
        RECT 399.000 182.000 399.500 182.500 ;
        RECT 400.500 181.750 401.500 185.000 ;
        RECT 397.000 181.250 401.500 181.750 ;
        RECT 397.000 178.000 398.000 181.250 ;
        RECT 398.250 180.000 398.750 180.500 ;
        RECT 399.000 180.250 399.500 180.750 ;
        RECT 399.750 180.000 400.250 180.500 ;
        RECT 398.250 179.000 398.790 180.000 ;
        RECT 399.000 179.000 399.500 180.000 ;
        RECT 399.710 179.000 400.250 180.000 ;
        RECT 399.000 178.250 399.500 178.750 ;
        RECT 400.500 178.000 401.500 181.250 ;
        RECT 397.000 177.500 401.500 178.000 ;
        RECT 397.000 174.250 398.000 177.500 ;
        RECT 398.250 176.250 398.750 176.750 ;
        RECT 399.000 176.500 399.500 177.000 ;
        RECT 399.750 176.250 400.250 176.750 ;
        RECT 398.250 175.250 398.790 176.250 ;
        RECT 399.000 175.250 399.500 176.250 ;
        RECT 399.710 175.250 400.250 176.250 ;
        RECT 399.000 174.500 399.500 175.000 ;
        RECT 400.500 174.250 401.500 177.500 ;
        RECT 397.000 173.750 401.500 174.250 ;
        RECT 397.000 170.500 398.000 173.750 ;
        RECT 398.250 172.500 398.750 173.000 ;
        RECT 399.000 172.750 399.500 173.250 ;
        RECT 399.750 172.500 400.250 173.000 ;
        RECT 398.250 171.500 398.790 172.500 ;
        RECT 399.000 171.500 399.500 172.500 ;
        RECT 399.710 171.500 400.250 172.500 ;
        RECT 399.000 170.750 399.500 171.250 ;
        RECT 400.500 170.500 401.500 173.750 ;
        RECT 397.000 170.000 401.500 170.500 ;
        RECT 397.000 166.750 398.000 170.000 ;
        RECT 398.250 168.750 398.750 169.250 ;
        RECT 399.000 169.000 399.500 169.500 ;
        RECT 399.750 168.750 400.250 169.250 ;
        RECT 398.250 167.750 398.790 168.750 ;
        RECT 399.000 167.750 399.500 168.750 ;
        RECT 399.710 167.750 400.250 168.750 ;
        RECT 399.000 167.000 399.500 167.500 ;
        RECT 400.500 166.750 401.500 170.000 ;
        RECT 397.000 166.250 401.500 166.750 ;
        RECT 406.500 193.000 407.500 196.000 ;
        RECT 407.750 195.000 408.250 195.500 ;
        RECT 408.500 195.250 409.000 195.750 ;
        RECT 409.250 195.000 409.750 195.500 ;
        RECT 407.750 194.000 408.290 195.000 ;
        RECT 408.500 194.000 409.000 195.000 ;
        RECT 409.210 194.000 409.750 195.000 ;
        RECT 408.500 193.250 409.000 193.750 ;
        RECT 410.000 193.000 411.000 196.000 ;
        RECT 406.500 192.500 411.000 193.000 ;
        RECT 406.500 189.250 407.500 192.500 ;
        RECT 407.750 191.250 408.250 191.750 ;
        RECT 408.500 191.500 409.000 192.000 ;
        RECT 409.250 191.250 409.750 191.750 ;
        RECT 407.750 190.250 408.290 191.250 ;
        RECT 408.500 190.250 409.000 191.250 ;
        RECT 409.210 190.250 409.750 191.250 ;
        RECT 408.500 189.500 409.000 190.000 ;
        RECT 410.000 189.250 411.000 192.500 ;
        RECT 406.500 188.750 411.000 189.250 ;
        RECT 406.500 185.500 407.500 188.750 ;
        RECT 407.750 187.500 408.250 188.000 ;
        RECT 408.500 187.750 409.000 188.250 ;
        RECT 409.250 187.500 409.750 188.000 ;
        RECT 407.750 186.500 408.290 187.500 ;
        RECT 408.500 186.500 409.000 187.500 ;
        RECT 409.210 186.500 409.750 187.500 ;
        RECT 408.500 185.750 409.000 186.250 ;
        RECT 410.000 185.500 411.000 188.750 ;
        RECT 406.500 185.000 411.000 185.500 ;
        RECT 406.500 181.750 407.500 185.000 ;
        RECT 407.750 183.750 408.250 184.250 ;
        RECT 408.500 184.000 409.000 184.500 ;
        RECT 409.250 183.750 409.750 184.250 ;
        RECT 407.750 182.750 408.290 183.750 ;
        RECT 408.500 182.750 409.000 183.750 ;
        RECT 409.210 182.750 409.750 183.750 ;
        RECT 408.500 182.000 409.000 182.500 ;
        RECT 410.000 181.750 411.000 185.000 ;
        RECT 406.500 181.250 411.000 181.750 ;
        RECT 406.500 178.000 407.500 181.250 ;
        RECT 407.750 180.000 408.250 180.500 ;
        RECT 408.500 180.250 409.000 180.750 ;
        RECT 409.250 180.000 409.750 180.500 ;
        RECT 407.750 179.000 408.290 180.000 ;
        RECT 408.500 179.000 409.000 180.000 ;
        RECT 409.210 179.000 409.750 180.000 ;
        RECT 408.500 178.250 409.000 178.750 ;
        RECT 410.000 178.000 411.000 181.250 ;
        RECT 406.500 177.500 411.000 178.000 ;
        RECT 406.500 174.250 407.500 177.500 ;
        RECT 407.750 176.250 408.250 176.750 ;
        RECT 408.500 176.500 409.000 177.000 ;
        RECT 409.250 176.250 409.750 176.750 ;
        RECT 407.750 175.250 408.290 176.250 ;
        RECT 408.500 175.250 409.000 176.250 ;
        RECT 409.210 175.250 409.750 176.250 ;
        RECT 408.500 174.500 409.000 175.000 ;
        RECT 410.000 174.250 411.000 177.500 ;
        RECT 406.500 173.750 411.000 174.250 ;
        RECT 406.500 170.500 407.500 173.750 ;
        RECT 407.750 172.500 408.250 173.000 ;
        RECT 408.500 172.750 409.000 173.250 ;
        RECT 409.250 172.500 409.750 173.000 ;
        RECT 407.750 171.500 408.290 172.500 ;
        RECT 408.500 171.500 409.000 172.500 ;
        RECT 409.210 171.500 409.750 172.500 ;
        RECT 408.500 170.750 409.000 171.250 ;
        RECT 410.000 170.500 411.000 173.750 ;
        RECT 406.500 170.000 411.000 170.500 ;
        RECT 406.500 166.750 407.500 170.000 ;
        RECT 407.750 168.750 408.250 169.250 ;
        RECT 408.500 169.000 409.000 169.500 ;
        RECT 409.250 168.750 409.750 169.250 ;
        RECT 407.750 167.750 408.290 168.750 ;
        RECT 408.500 167.750 409.000 168.750 ;
        RECT 409.210 167.750 409.750 168.750 ;
        RECT 408.500 167.000 409.000 167.500 ;
        RECT 410.000 166.750 411.000 170.000 ;
        RECT 406.500 166.250 411.000 166.750 ;
        RECT 301.920 165.780 312.640 165.920 ;
        RECT 297.230 165.720 297.550 165.780 ;
        RECT 297.705 165.735 297.995 165.780 ;
        RECT 301.415 165.720 301.735 165.780 ;
        RECT 300.450 165.380 300.770 165.640 ;
        RECT 311.965 165.580 312.255 165.625 ;
        RECT 301.920 165.440 312.255 165.580 ;
        RECT 298.610 165.040 298.930 165.300 ;
        RECT 299.530 165.240 299.850 165.300 ;
        RECT 301.920 165.285 302.060 165.440 ;
        RECT 311.965 165.395 312.255 165.440 ;
        RECT 301.845 165.240 302.135 165.285 ;
        RECT 299.530 165.100 302.135 165.240 ;
        RECT 299.530 165.040 299.850 165.100 ;
        RECT 301.845 165.055 302.135 165.100 ;
        RECT 302.765 165.055 303.055 165.285 ;
        RECT 310.585 165.240 310.875 165.285 ;
        RECT 311.490 165.240 311.810 165.300 ;
        RECT 312.500 165.240 312.640 165.780 ;
        RECT 310.585 165.100 312.640 165.240 ;
        RECT 310.585 165.055 310.875 165.100 ;
        RECT 298.150 164.900 298.470 164.960 ;
        RECT 302.840 164.900 302.980 165.055 ;
        RECT 311.490 165.040 311.810 165.100 ;
        RECT 379.000 165.000 411.250 166.000 ;
        RECT 311.045 164.900 311.335 164.945 ;
        RECT 298.150 164.760 311.335 164.900 ;
        RECT 298.150 164.700 298.470 164.760 ;
        RECT 311.045 164.715 311.335 164.760 ;
        RECT 291.500 164.080 320.500 164.560 ;
        RECT 298.150 163.680 298.470 163.940 ;
        RECT 311.490 163.880 311.810 163.940 ;
        RECT 311.965 163.880 312.255 163.925 ;
        RECT 311.490 163.740 312.255 163.880 ;
        RECT 311.490 163.680 311.810 163.740 ;
        RECT 311.965 163.695 312.255 163.740 ;
        RECT 296.770 163.540 297.090 163.600 ;
        RECT 298.625 163.540 298.915 163.585 ;
        RECT 296.770 163.400 301.140 163.540 ;
        RECT 296.770 163.340 297.090 163.400 ;
        RECT 298.625 163.355 298.915 163.400 ;
        RECT 297.230 163.000 297.550 163.260 ;
        RECT 300.450 163.000 300.770 163.260 ;
        RECT 301.000 163.245 301.140 163.400 ;
        RECT 379.250 163.500 390.250 164.000 ;
        RECT 300.925 163.200 301.215 163.245 ;
        RECT 310.570 163.200 310.890 163.260 ;
        RECT 311.505 163.200 311.795 163.245 ;
        RECT 300.925 163.060 311.795 163.200 ;
        RECT 300.925 163.015 301.215 163.060 ;
        RECT 310.570 163.000 310.890 163.060 ;
        RECT 311.505 163.015 311.795 163.060 ;
        RECT 312.885 163.200 313.175 163.245 ;
        RECT 314.250 163.200 314.570 163.260 ;
        RECT 312.885 163.060 314.570 163.200 ;
        RECT 312.885 163.015 313.175 163.060 ;
        RECT 314.250 163.000 314.570 163.060 ;
        RECT 299.530 162.320 299.850 162.580 ;
        RECT 313.790 162.320 314.110 162.580 ;
        RECT 294.470 161.980 294.790 162.240 ;
        RECT 296.310 162.180 296.630 162.240 ;
        RECT 300.940 162.180 301.260 162.240 ;
        RECT 296.310 162.040 301.260 162.180 ;
        RECT 296.310 161.980 296.630 162.040 ;
        RECT 300.940 161.980 301.260 162.040 ;
        RECT 290.000 161.360 320.500 161.840 ;
        RECT 291.500 158.640 320.500 159.120 ;
        RECT 299.250 156.000 378.000 158.000 ;
        RECT 285.500 153.500 354.750 155.500 ;
        RECT 379.250 153.000 379.750 163.500 ;
        RECT 380.750 162.750 381.750 163.250 ;
        RECT 380.000 154.000 380.720 162.500 ;
        RECT 381.780 154.000 382.500 162.500 ;
        RECT 380.750 153.250 381.750 153.750 ;
        RECT 382.750 153.000 383.250 163.500 ;
        RECT 384.250 162.750 385.250 163.250 ;
        RECT 383.500 154.000 384.220 162.500 ;
        RECT 385.280 154.000 386.000 162.500 ;
        RECT 384.250 153.250 385.250 153.750 ;
        RECT 386.250 153.000 386.750 163.500 ;
        RECT 387.750 162.750 388.750 163.250 ;
        RECT 387.000 154.000 387.720 162.500 ;
        RECT 388.780 154.000 389.500 162.500 ;
        RECT 389.750 158.000 390.250 163.500 ;
        RECT 390.750 159.000 391.250 165.000 ;
        RECT 391.585 160.750 391.815 165.000 ;
        RECT 392.045 160.500 392.275 164.750 ;
        RECT 392.505 160.750 392.735 165.000 ;
        RECT 392.965 160.500 393.195 164.750 ;
        RECT 393.425 160.750 393.655 165.000 ;
        RECT 393.885 160.500 394.115 164.750 ;
        RECT 394.345 160.750 394.575 165.000 ;
        RECT 394.805 160.500 395.035 164.750 ;
        RECT 395.265 160.750 395.495 165.000 ;
        RECT 395.725 160.500 395.955 164.750 ;
        RECT 396.185 160.750 396.415 165.000 ;
        RECT 392.045 160.000 395.955 160.500 ;
        RECT 393.750 159.250 394.250 159.750 ;
        RECT 396.750 159.000 397.250 165.000 ;
        RECT 397.585 160.750 397.815 165.000 ;
        RECT 398.045 160.500 398.275 164.750 ;
        RECT 398.505 160.750 398.735 165.000 ;
        RECT 398.965 160.500 399.195 164.750 ;
        RECT 399.425 160.750 399.655 165.000 ;
        RECT 399.885 160.500 400.115 164.750 ;
        RECT 400.345 160.750 400.575 165.000 ;
        RECT 400.805 160.500 401.035 164.750 ;
        RECT 401.265 160.750 401.495 165.000 ;
        RECT 401.725 160.500 401.955 164.750 ;
        RECT 402.185 160.750 402.415 165.000 ;
        RECT 398.045 160.000 401.955 160.500 ;
        RECT 399.750 159.250 400.250 159.750 ;
        RECT 402.750 159.000 403.250 165.000 ;
        RECT 403.585 160.750 403.815 165.000 ;
        RECT 404.045 160.500 404.275 164.750 ;
        RECT 404.505 160.750 404.735 165.000 ;
        RECT 404.965 160.500 405.195 164.750 ;
        RECT 405.425 160.750 405.655 165.000 ;
        RECT 405.885 160.500 406.115 164.750 ;
        RECT 406.345 160.750 406.575 165.000 ;
        RECT 406.805 160.500 407.035 164.750 ;
        RECT 407.265 160.750 407.495 165.000 ;
        RECT 407.725 160.500 407.955 164.750 ;
        RECT 408.185 160.750 408.415 165.000 ;
        RECT 408.750 164.000 409.750 165.000 ;
        RECT 408.750 163.000 421.000 164.000 ;
        RECT 404.045 160.000 407.955 160.500 ;
        RECT 405.750 159.250 406.250 159.750 ;
        RECT 408.750 159.000 409.250 163.000 ;
        RECT 390.750 158.500 409.250 159.000 ;
        RECT 409.500 159.000 410.000 163.000 ;
        RECT 410.185 160.750 410.415 163.000 ;
        RECT 410.625 160.500 410.855 162.750 ;
        RECT 411.065 160.750 411.295 163.000 ;
        RECT 411.505 160.500 411.735 162.750 ;
        RECT 411.945 160.750 412.175 163.000 ;
        RECT 412.385 160.500 412.615 162.750 ;
        RECT 412.825 160.750 413.055 163.000 ;
        RECT 413.265 160.500 413.495 162.750 ;
        RECT 413.705 160.750 413.935 163.000 ;
        RECT 414.145 160.500 414.375 162.750 ;
        RECT 414.585 160.750 414.815 163.000 ;
        RECT 410.625 160.000 414.375 160.500 ;
        RECT 412.250 159.250 412.750 159.750 ;
        RECT 415.000 159.000 415.500 163.000 ;
        RECT 415.685 160.750 415.915 163.000 ;
        RECT 416.125 160.500 416.355 162.750 ;
        RECT 416.565 160.750 416.795 163.000 ;
        RECT 417.005 160.500 417.235 162.750 ;
        RECT 417.445 160.750 417.675 163.000 ;
        RECT 417.885 160.500 418.115 162.750 ;
        RECT 418.325 160.750 418.555 163.000 ;
        RECT 418.765 160.500 418.995 162.750 ;
        RECT 419.205 160.750 419.435 163.000 ;
        RECT 419.645 160.500 419.875 162.750 ;
        RECT 420.085 160.750 420.315 163.000 ;
        RECT 416.125 160.000 419.875 160.500 ;
        RECT 417.750 159.250 418.250 159.750 ;
        RECT 420.500 159.000 421.000 163.000 ;
        RECT 409.500 158.500 421.000 159.000 ;
        RECT 389.750 157.500 409.250 158.000 ;
        RECT 387.750 153.250 388.750 153.750 ;
        RECT 389.750 153.000 391.250 157.500 ;
        RECT 393.750 156.750 394.250 157.250 ;
        RECT 392.045 156.000 395.955 156.500 ;
        RECT 285.500 151.000 354.750 153.000 ;
        RECT 379.250 152.500 391.250 153.000 ;
        RECT 379.250 151.500 379.750 152.500 ;
        RECT 382.750 151.500 383.250 152.500 ;
        RECT 386.250 151.500 386.750 152.500 ;
        RECT 389.750 151.500 391.250 152.500 ;
        RECT 391.585 151.500 391.815 155.750 ;
        RECT 392.045 151.750 392.275 156.000 ;
        RECT 392.505 151.500 392.735 155.750 ;
        RECT 392.965 151.750 393.195 156.000 ;
        RECT 393.425 151.500 393.655 155.750 ;
        RECT 393.885 151.750 394.115 156.000 ;
        RECT 394.345 151.500 394.575 155.750 ;
        RECT 394.805 151.750 395.035 156.000 ;
        RECT 395.265 151.500 395.495 155.750 ;
        RECT 395.725 151.750 395.955 156.000 ;
        RECT 396.185 151.500 396.415 155.750 ;
        RECT 396.750 151.500 397.250 157.500 ;
        RECT 399.750 156.750 400.250 157.250 ;
        RECT 398.045 156.000 401.955 156.500 ;
        RECT 397.585 151.500 397.815 155.750 ;
        RECT 398.045 151.750 398.275 156.000 ;
        RECT 398.505 151.500 398.735 155.750 ;
        RECT 398.965 151.750 399.195 156.000 ;
        RECT 399.425 151.500 399.655 155.750 ;
        RECT 399.885 151.750 400.115 156.000 ;
        RECT 400.345 151.500 400.575 155.750 ;
        RECT 400.805 151.750 401.035 156.000 ;
        RECT 401.265 151.500 401.495 155.750 ;
        RECT 401.725 151.750 401.955 156.000 ;
        RECT 402.185 151.500 402.415 155.750 ;
        RECT 402.750 151.500 403.250 157.500 ;
        RECT 405.750 156.750 406.250 157.250 ;
        RECT 404.045 156.000 407.955 156.500 ;
        RECT 403.585 151.500 403.815 155.750 ;
        RECT 404.045 151.750 404.275 156.000 ;
        RECT 404.505 151.500 404.735 155.750 ;
        RECT 404.965 151.750 405.195 156.000 ;
        RECT 405.425 151.500 405.655 155.750 ;
        RECT 405.885 151.750 406.115 156.000 ;
        RECT 406.345 151.500 406.575 155.750 ;
        RECT 406.805 151.750 407.035 156.000 ;
        RECT 407.265 151.500 407.495 155.750 ;
        RECT 407.725 151.750 407.955 156.000 ;
        RECT 408.185 151.500 408.415 155.750 ;
        RECT 408.750 153.500 409.250 157.500 ;
        RECT 409.500 157.500 421.000 158.000 ;
        RECT 409.500 153.500 410.000 157.500 ;
        RECT 412.250 156.750 412.750 157.250 ;
        RECT 410.625 156.000 414.375 156.500 ;
        RECT 410.185 153.500 410.415 155.825 ;
        RECT 410.625 153.825 410.855 156.000 ;
        RECT 411.065 153.500 411.295 155.825 ;
        RECT 411.505 153.825 411.735 156.000 ;
        RECT 411.945 153.500 412.175 155.825 ;
        RECT 412.385 153.825 412.615 156.000 ;
        RECT 412.825 153.500 413.055 155.825 ;
        RECT 413.265 153.825 413.495 156.000 ;
        RECT 413.705 153.500 413.935 155.825 ;
        RECT 414.145 153.825 414.375 156.000 ;
        RECT 414.585 153.500 414.815 155.825 ;
        RECT 415.000 153.500 415.500 157.500 ;
        RECT 417.750 156.750 418.250 157.250 ;
        RECT 416.125 156.000 419.875 156.500 ;
        RECT 415.685 153.500 415.915 155.825 ;
        RECT 416.125 153.825 416.355 156.000 ;
        RECT 416.565 153.500 416.795 155.825 ;
        RECT 417.005 153.825 417.235 156.000 ;
        RECT 417.445 153.500 417.675 155.825 ;
        RECT 417.885 153.825 418.115 156.000 ;
        RECT 418.325 153.500 418.555 155.825 ;
        RECT 418.765 153.825 418.995 156.000 ;
        RECT 419.205 153.500 419.435 155.825 ;
        RECT 419.645 153.825 419.875 156.000 ;
        RECT 420.085 153.500 420.315 155.825 ;
        RECT 420.500 153.500 421.000 157.500 ;
        RECT 408.750 152.500 421.000 153.500 ;
        RECT 408.750 151.500 409.750 152.500 ;
        RECT 286.000 144.500 287.000 151.000 ;
        RECT 289.500 149.500 301.250 150.750 ;
        RECT 307.750 150.250 339.500 150.750 ;
        RECT 311.500 149.500 340.250 150.000 ;
        RECT 296.000 148.750 304.250 149.250 ;
        RECT 310.750 148.750 319.500 149.250 ;
        RECT 287.250 148.000 353.500 148.500 ;
        RECT 287.970 147.750 290.160 147.830 ;
        RECT 287.970 147.600 290.750 147.750 ;
        RECT 292.970 147.600 295.160 147.830 ;
        RECT 303.970 147.600 306.160 147.830 ;
        RECT 308.970 147.750 311.160 147.830 ;
        RECT 317.220 147.750 319.410 147.830 ;
        RECT 308.970 147.600 311.250 147.750 ;
        RECT 317.220 147.600 319.500 147.750 ;
        RECT 324.720 147.600 326.910 147.830 ;
        RECT 329.720 147.600 331.910 147.830 ;
        RECT 335.470 147.600 337.660 147.830 ;
        RECT 289.500 147.000 290.750 147.600 ;
        RECT 291.750 147.395 292.250 147.500 ;
        RECT 287.750 146.500 290.750 147.000 ;
        RECT 291.740 147.250 292.250 147.395 ;
        RECT 294.500 147.250 295.000 147.600 ;
        RECT 291.740 147.000 295.000 147.250 ;
        RECT 291.740 146.500 296.500 147.000 ;
        RECT 288.310 145.905 291.600 146.135 ;
        RECT 291.300 145.095 291.530 145.545 ;
        RECT 291.740 145.095 292.250 146.500 ;
        RECT 293.250 145.750 294.250 146.250 ;
        RECT 291.750 145.000 292.250 145.095 ;
        RECT 294.500 144.915 295.000 146.500 ;
        RECT 296.740 146.250 296.970 147.395 ;
        RECT 298.525 146.750 298.980 147.395 ;
        RECT 300.660 146.750 300.890 147.395 ;
        RECT 303.160 146.750 303.390 147.395 ;
        RECT 305.500 147.000 306.000 147.600 ;
        RECT 298.525 146.495 300.250 146.750 ;
        RECT 298.750 146.250 300.250 146.495 ;
        RECT 296.740 145.750 298.500 146.250 ;
        RECT 298.750 145.750 299.250 146.250 ;
        RECT 299.750 146.105 300.250 146.250 ;
        RECT 300.500 146.250 301.750 146.750 ;
        RECT 300.500 146.105 301.000 146.250 ;
        RECT 296.300 145.095 296.530 145.545 ;
        RECT 296.740 145.095 296.970 145.750 ;
        RECT 298.750 145.545 298.980 145.750 ;
        RECT 298.525 145.095 298.980 145.545 ;
        RECT 299.750 145.705 300.900 145.935 ;
        RECT 301.250 145.750 301.750 146.250 ;
        RECT 302.250 146.105 302.750 146.750 ;
        RECT 303.000 146.305 303.500 146.750 ;
        RECT 303.750 146.500 306.000 147.000 ;
        RECT 303.000 146.075 304.750 146.305 ;
        RECT 302.250 145.750 303.400 145.935 ;
        RECT 304.250 145.750 304.750 146.075 ;
        RECT 301.250 145.705 303.400 145.750 ;
        RECT 299.750 145.250 300.250 145.705 ;
        RECT 301.250 145.250 302.750 145.705 ;
        RECT 305.500 144.915 306.000 146.500 ;
        RECT 307.740 147.000 307.970 147.395 ;
        RECT 310.750 147.000 311.250 147.600 ;
        RECT 307.740 146.500 311.250 147.000 ;
        RECT 307.740 145.750 308.250 146.500 ;
        RECT 309.250 145.750 310.500 146.250 ;
        RECT 307.300 145.095 307.530 145.545 ;
        RECT 307.740 145.095 307.970 145.750 ;
        RECT 310.750 144.915 311.250 146.500 ;
        RECT 312.740 146.250 312.970 147.395 ;
        RECT 312.740 145.750 313.250 146.250 ;
        RECT 314.750 146.090 315.250 146.750 ;
        RECT 315.390 146.295 315.620 147.395 ;
        RECT 315.390 146.065 315.860 146.295 ;
        RECT 316.170 146.250 316.400 147.395 ;
        RECT 319.000 147.000 319.500 147.600 ;
        RECT 343.000 147.395 345.250 147.500 ;
        RECT 317.340 146.500 319.500 147.000 ;
        RECT 314.750 145.750 315.250 145.935 ;
        RECT 312.300 145.095 312.530 145.545 ;
        RECT 312.740 145.250 315.250 145.750 ;
        RECT 312.740 145.095 312.970 145.250 ;
        RECT 315.390 145.095 315.620 146.065 ;
        RECT 316.000 145.750 318.000 146.250 ;
        RECT 316.170 145.095 316.400 145.750 ;
        RECT 319.000 144.915 319.500 146.500 ;
        RECT 320.990 146.250 321.220 147.395 ;
        RECT 322.775 147.000 323.230 147.395 ;
        RECT 328.490 147.000 328.720 147.395 ;
        RECT 333.490 147.000 333.720 147.395 ;
        RECT 339.240 147.000 339.470 147.395 ;
        RECT 322.775 146.500 325.500 147.000 ;
        RECT 328.490 146.500 330.500 147.000 ;
        RECT 333.490 146.500 336.250 147.000 ;
        RECT 322.775 146.495 323.500 146.500 ;
        RECT 320.990 145.750 322.750 146.250 ;
        RECT 323.000 145.750 323.500 146.495 ;
        RECT 325.060 145.905 328.350 146.135 ;
        RECT 328.490 145.750 329.000 146.500 ;
        RECT 330.060 145.905 333.350 146.135 ;
        RECT 333.490 145.750 334.000 146.500 ;
        RECT 339.240 146.250 340.750 147.000 ;
        RECT 341.025 146.495 341.480 147.395 ;
        RECT 342.775 146.495 345.250 147.395 ;
        RECT 341.250 146.250 341.480 146.495 ;
        RECT 335.810 145.905 339.100 146.135 ;
        RECT 339.240 145.750 341.000 146.250 ;
        RECT 341.250 145.750 342.750 146.250 ;
        RECT 320.550 145.095 320.780 145.545 ;
        RECT 320.990 145.095 321.220 145.750 ;
        RECT 323.000 145.545 323.230 145.750 ;
        RECT 322.775 145.095 323.230 145.545 ;
        RECT 328.050 145.095 328.280 145.545 ;
        RECT 328.490 145.095 328.720 145.750 ;
        RECT 333.050 145.095 333.280 145.545 ;
        RECT 333.490 145.095 333.720 145.750 ;
        RECT 338.800 145.095 339.030 145.545 ;
        RECT 339.240 145.095 339.470 145.750 ;
        RECT 341.250 145.545 341.480 145.750 ;
        RECT 343.000 145.545 345.250 146.495 ;
        RECT 341.025 145.095 341.480 145.545 ;
        RECT 342.775 145.095 345.250 145.545 ;
        RECT 343.000 145.000 345.250 145.095 ;
        RECT 287.970 144.685 290.880 144.915 ;
        RECT 292.970 144.685 295.880 144.915 ;
        RECT 303.970 144.685 306.880 144.915 ;
        RECT 308.970 144.685 311.880 144.915 ;
        RECT 317.220 144.685 320.130 144.915 ;
        RECT 324.720 144.685 327.630 144.915 ;
        RECT 329.720 144.685 332.630 144.915 ;
        RECT 335.470 144.685 338.380 144.915 ;
        RECT 353.750 144.500 354.750 151.000 ;
        RECT 379.000 150.500 411.250 151.500 ;
        RECT 359.500 149.750 381.750 150.250 ;
        RECT 387.500 149.750 392.000 150.500 ;
        RECT 387.500 146.500 388.500 149.750 ;
        RECT 389.500 149.000 390.000 149.500 ;
        RECT 388.750 147.750 389.290 148.750 ;
        RECT 389.500 147.750 390.000 148.750 ;
        RECT 390.210 147.750 390.750 148.750 ;
        RECT 388.750 147.250 389.250 147.750 ;
        RECT 389.500 147.000 390.000 147.500 ;
        RECT 390.250 147.250 390.750 147.750 ;
        RECT 391.000 146.500 392.000 149.750 ;
        RECT 361.500 146.000 381.750 146.500 ;
        RECT 387.500 146.000 392.000 146.500 ;
        RECT 286.000 144.000 354.750 144.500 ;
        RECT 286.000 137.500 287.000 144.000 ;
        RECT 293.750 143.250 308.250 143.750 ;
        RECT 310.000 143.250 323.500 143.750 ;
        RECT 294.000 142.500 300.250 143.000 ;
        RECT 314.000 142.500 340.250 143.000 ;
        RECT 314.750 141.750 329.000 142.250 ;
        RECT 292.250 141.000 353.500 141.500 ;
        RECT 300.500 140.535 308.000 140.765 ;
        RECT 315.750 140.750 317.860 140.860 ;
        RECT 294.270 139.495 294.725 140.395 ;
        RECT 296.020 139.495 296.400 140.395 ;
        RECT 296.540 139.890 297.710 140.120 ;
        RECT 294.270 139.250 294.500 139.495 ;
        RECT 296.020 139.250 296.250 139.495 ;
        RECT 296.540 139.290 296.770 139.890 ;
        RECT 294.000 138.750 294.500 139.250 ;
        RECT 294.750 138.750 295.500 139.250 ;
        RECT 295.750 138.750 296.250 139.250 ;
        RECT 296.390 138.975 296.770 139.290 ;
        RECT 297.250 139.250 299.000 139.750 ;
        RECT 299.350 139.250 299.580 140.395 ;
        RECT 300.130 139.295 300.360 140.395 ;
        RECT 297.250 139.105 297.750 139.250 ;
        RECT 294.270 138.545 294.500 138.750 ;
        RECT 296.020 138.545 296.250 138.750 ;
        RECT 294.270 138.095 294.725 138.545 ;
        RECT 296.020 138.095 296.400 138.545 ;
        RECT 296.540 138.110 296.770 138.975 ;
        RECT 297.250 138.750 297.750 138.935 ;
        RECT 299.250 138.750 299.750 139.250 ;
        RECT 299.890 139.065 300.360 139.295 ;
        RECT 300.500 139.090 301.000 140.535 ;
        RECT 307.500 140.395 308.000 140.535 ;
        RECT 315.500 140.630 317.860 140.750 ;
        RECT 301.770 139.495 302.225 140.395 ;
        RECT 304.270 139.495 304.725 140.395 ;
        RECT 306.020 139.495 306.475 140.395 ;
        RECT 307.500 139.495 308.225 140.395 ;
        RECT 309.520 139.495 309.975 140.395 ;
        RECT 315.500 140.250 316.250 140.630 ;
        RECT 316.840 140.200 317.070 140.630 ;
        RECT 318.480 140.000 318.710 140.860 ;
        RECT 323.895 140.630 325.015 140.860 ;
        RECT 325.465 140.630 326.765 140.860 ;
        RECT 328.750 140.750 330.860 140.860 ;
        RECT 315.600 139.770 318.710 140.000 ;
        RECT 315.600 139.500 317.000 139.770 ;
        RECT 301.770 139.250 302.000 139.495 ;
        RECT 304.270 139.250 304.500 139.495 ;
        RECT 306.020 139.250 306.250 139.495 ;
        RECT 307.500 139.250 308.000 139.495 ;
        RECT 309.520 139.250 309.750 139.495 ;
        RECT 297.250 138.250 299.580 138.750 ;
        RECT 296.540 137.880 297.310 138.110 ;
        RECT 299.350 138.095 299.580 138.250 ;
        RECT 300.130 138.095 300.360 139.065 ;
        RECT 300.500 138.750 301.000 138.935 ;
        RECT 301.500 138.750 302.000 139.250 ;
        RECT 302.250 138.750 304.500 139.250 ;
        RECT 304.750 138.750 306.250 139.250 ;
        RECT 306.500 138.750 308.000 139.250 ;
        RECT 308.250 138.750 309.750 139.250 ;
        RECT 310.000 138.750 312.000 139.250 ;
        RECT 315.750 138.750 316.250 139.250 ;
        RECT 317.250 138.920 317.480 139.320 ;
        RECT 317.690 139.060 319.360 139.290 ;
        RECT 319.500 139.250 319.730 140.395 ;
        RECT 322.025 139.495 322.480 140.395 ;
        RECT 322.250 139.335 322.480 139.495 ;
        RECT 323.250 139.335 323.750 139.750 ;
        RECT 323.895 139.495 324.125 140.630 ;
        RECT 324.745 140.260 325.915 140.490 ;
        RECT 325.185 139.660 326.395 140.120 ;
        RECT 325.935 139.335 326.395 139.660 ;
        RECT 326.535 139.495 326.765 140.630 ;
        RECT 328.500 140.630 330.860 140.750 ;
        RECT 328.500 140.250 329.250 140.630 ;
        RECT 329.840 140.200 330.070 140.630 ;
        RECT 331.480 140.000 331.710 140.860 ;
        RECT 336.895 140.630 338.015 140.860 ;
        RECT 338.465 140.630 339.765 140.860 ;
        RECT 328.600 139.770 331.710 140.000 ;
        RECT 328.600 139.500 330.000 139.770 ;
        RECT 319.500 139.020 322.000 139.250 ;
        RECT 322.230 139.105 325.045 139.335 ;
        RECT 300.500 138.545 302.000 138.750 ;
        RECT 304.270 138.545 304.500 138.750 ;
        RECT 306.020 138.545 306.250 138.750 ;
        RECT 307.770 138.545 308.000 138.750 ;
        RECT 309.520 138.545 309.750 138.750 ;
        RECT 317.250 138.690 318.480 138.920 ;
        RECT 319.500 138.750 320.000 139.020 ;
        RECT 321.500 138.750 322.000 139.020 ;
        RECT 322.250 138.750 322.750 139.105 ;
        RECT 325.250 138.965 325.750 139.250 ;
        RECT 325.935 139.105 327.250 139.335 ;
        RECT 300.500 138.250 302.225 138.545 ;
        RECT 301.770 138.095 302.225 138.250 ;
        RECT 304.270 138.095 304.725 138.545 ;
        RECT 306.020 138.095 306.475 138.545 ;
        RECT 307.770 138.095 308.225 138.545 ;
        RECT 309.520 138.095 309.975 138.545 ;
        RECT 315.980 138.315 317.020 138.545 ;
        RECT 317.260 138.315 318.980 138.545 ;
        RECT 315.980 138.095 316.210 138.315 ;
        RECT 317.260 138.095 317.490 138.315 ;
        RECT 319.500 138.095 319.730 138.750 ;
        RECT 322.250 138.545 322.480 138.750 ;
        RECT 322.025 138.095 322.480 138.545 ;
        RECT 323.250 138.735 326.415 138.965 ;
        RECT 326.750 138.750 327.250 139.105 ;
        RECT 328.750 138.750 329.250 139.250 ;
        RECT 330.250 138.920 330.480 139.320 ;
        RECT 330.690 139.060 332.360 139.290 ;
        RECT 332.500 139.250 332.730 140.395 ;
        RECT 335.025 139.495 335.480 140.395 ;
        RECT 335.250 139.335 335.480 139.495 ;
        RECT 336.250 139.335 336.750 139.750 ;
        RECT 336.895 139.495 337.125 140.630 ;
        RECT 337.745 140.260 338.915 140.490 ;
        RECT 338.185 139.660 339.395 140.120 ;
        RECT 338.935 139.335 339.395 139.660 ;
        RECT 339.535 139.495 339.765 140.630 ;
        RECT 348.250 140.395 349.250 140.500 ;
        RECT 332.500 139.020 335.000 139.250 ;
        RECT 335.230 139.105 338.045 139.335 ;
        RECT 323.250 138.250 323.750 138.735 ;
        RECT 330.250 138.690 331.480 138.920 ;
        RECT 332.500 138.750 333.000 139.020 ;
        RECT 334.500 138.750 335.000 139.020 ;
        RECT 335.250 138.750 335.750 139.105 ;
        RECT 338.250 138.965 338.750 139.250 ;
        RECT 338.935 139.105 340.250 139.335 ;
        RECT 342.250 139.250 344.250 139.750 ;
        RECT 344.400 139.495 344.980 140.395 ;
        RECT 346.025 139.495 346.480 140.395 ;
        RECT 347.525 139.495 347.980 140.395 ;
        RECT 348.250 139.500 350.480 140.395 ;
        RECT 350.025 139.495 350.480 139.500 ;
        RECT 323.935 137.870 324.165 138.545 ;
        RECT 326.495 138.240 326.725 138.545 ;
        RECT 324.845 138.010 326.725 138.240 ;
        RECT 328.980 138.315 330.020 138.545 ;
        RECT 330.260 138.315 331.980 138.545 ;
        RECT 328.980 138.095 329.210 138.315 ;
        RECT 330.260 138.095 330.490 138.315 ;
        RECT 332.500 138.095 332.730 138.750 ;
        RECT 335.250 138.545 335.480 138.750 ;
        RECT 335.025 138.095 335.480 138.545 ;
        RECT 336.250 138.735 339.415 138.965 ;
        RECT 339.750 138.750 340.250 139.105 ;
        RECT 343.750 139.075 344.250 139.250 ;
        RECT 344.750 139.250 344.980 139.495 ;
        RECT 346.250 139.250 346.480 139.495 ;
        RECT 347.750 139.250 347.980 139.495 ;
        RECT 350.250 139.250 350.480 139.495 ;
        RECT 343.750 138.750 344.400 138.935 ;
        RECT 344.750 138.750 346.000 139.250 ;
        RECT 346.250 138.750 347.500 139.250 ;
        RECT 347.750 138.750 350.000 139.250 ;
        RECT 350.250 138.750 350.750 139.250 ;
        RECT 336.250 138.250 336.750 138.735 ;
        RECT 336.935 137.870 337.165 138.545 ;
        RECT 339.495 138.240 339.725 138.545 ;
        RECT 343.750 138.250 344.500 138.750 ;
        RECT 337.845 138.010 339.725 138.240 ;
        RECT 344.750 138.095 345.030 138.750 ;
        RECT 346.250 138.545 346.480 138.750 ;
        RECT 347.750 138.545 347.980 138.750 ;
        RECT 350.250 138.545 350.480 138.750 ;
        RECT 346.025 138.095 346.480 138.545 ;
        RECT 347.525 138.095 347.980 138.545 ;
        RECT 350.025 138.095 350.480 138.545 ;
        RECT 315.600 137.640 318.900 137.870 ;
        RECT 323.935 137.640 325.675 137.870 ;
        RECT 328.600 137.640 331.900 137.870 ;
        RECT 336.935 137.640 338.675 137.870 ;
        RECT 353.750 137.500 354.750 144.000 ;
        RECT 387.500 142.750 388.500 146.000 ;
        RECT 389.500 145.250 390.000 145.750 ;
        RECT 388.750 144.000 389.290 145.000 ;
        RECT 389.500 144.000 390.000 145.000 ;
        RECT 390.210 144.000 390.750 145.000 ;
        RECT 388.750 143.500 389.250 144.000 ;
        RECT 389.500 143.250 390.000 143.750 ;
        RECT 390.250 143.500 390.750 144.000 ;
        RECT 391.000 142.750 392.000 146.000 ;
        RECT 363.500 142.250 381.750 142.750 ;
        RECT 387.500 142.250 392.000 142.750 ;
        RECT 387.500 139.000 388.500 142.250 ;
        RECT 389.500 141.500 390.000 142.000 ;
        RECT 388.750 140.250 389.290 141.250 ;
        RECT 389.500 140.250 390.000 141.250 ;
        RECT 390.210 140.250 390.750 141.250 ;
        RECT 388.750 139.750 389.250 140.250 ;
        RECT 389.500 139.500 390.000 140.000 ;
        RECT 390.250 139.750 390.750 140.250 ;
        RECT 391.000 139.000 392.000 142.250 ;
        RECT 365.500 138.500 381.750 139.000 ;
        RECT 387.500 138.500 392.000 139.000 ;
        RECT 286.000 137.000 354.750 137.500 ;
        RECT 286.000 130.500 287.000 137.000 ;
        RECT 294.000 136.250 315.250 136.750 ;
        RECT 315.750 136.250 323.750 136.750 ;
        RECT 328.750 136.250 336.750 136.750 ;
        RECT 344.000 136.250 349.000 136.750 ;
        RECT 297.750 135.500 308.000 136.000 ;
        RECT 319.500 135.500 330.000 136.000 ;
        RECT 332.500 135.500 335.000 136.000 ;
        RECT 297.000 134.750 309.250 135.250 ;
        RECT 315.000 134.750 327.250 135.250 ;
        RECT 327.500 134.750 341.000 135.250 ;
        RECT 342.250 134.750 343.500 135.250 ;
        RECT 343.750 134.750 348.250 135.250 ;
        RECT 292.250 134.000 353.500 134.500 ;
        RECT 294.270 132.250 294.500 133.395 ;
        RECT 295.290 133.000 295.520 133.860 ;
        RECT 296.140 133.630 298.250 133.860 ;
        RECT 296.930 133.250 298.250 133.630 ;
        RECT 300.500 133.535 308.000 133.765 ;
        RECT 296.930 133.200 297.160 133.250 ;
        RECT 295.290 132.770 298.400 133.000 ;
        RECT 295.750 132.500 298.400 132.770 ;
        RECT 293.500 131.750 294.500 132.250 ;
        RECT 294.640 132.060 296.310 132.290 ;
        RECT 296.520 131.920 296.750 132.320 ;
        RECT 299.350 132.250 299.580 133.395 ;
        RECT 300.130 132.295 300.360 133.395 ;
        RECT 294.270 131.095 294.500 131.750 ;
        RECT 295.520 131.690 296.750 131.920 ;
        RECT 297.750 131.750 298.250 132.250 ;
        RECT 298.500 131.750 299.750 132.250 ;
        RECT 299.890 132.065 300.360 132.295 ;
        RECT 300.500 132.090 301.000 133.535 ;
        RECT 307.500 133.395 308.000 133.535 ;
        RECT 312.980 133.630 313.340 133.860 ;
        RECT 313.890 133.750 314.500 133.860 ;
        RECT 301.770 132.495 302.225 133.395 ;
        RECT 304.270 132.495 304.725 133.395 ;
        RECT 306.020 132.495 306.475 133.395 ;
        RECT 307.500 132.495 308.225 133.395 ;
        RECT 309.520 132.495 309.975 133.395 ;
        RECT 301.770 132.250 302.000 132.495 ;
        RECT 304.270 132.250 304.500 132.495 ;
        RECT 306.020 132.250 306.250 132.495 ;
        RECT 307.500 132.250 308.000 132.495 ;
        RECT 309.520 132.250 309.750 132.495 ;
        RECT 312.180 132.250 312.410 133.395 ;
        RECT 312.980 133.000 313.210 133.630 ;
        RECT 313.890 133.250 316.250 133.750 ;
        RECT 316.735 133.630 318.035 133.860 ;
        RECT 318.485 133.630 319.605 133.860 ;
        RECT 312.980 132.770 316.500 133.000 ;
        RECT 295.020 131.315 296.740 131.545 ;
        RECT 296.980 131.315 298.020 131.545 ;
        RECT 296.510 131.095 296.740 131.315 ;
        RECT 297.790 131.095 298.020 131.315 ;
        RECT 299.350 131.095 299.580 131.750 ;
        RECT 300.130 131.095 300.360 132.065 ;
        RECT 300.500 131.750 301.000 131.935 ;
        RECT 301.500 131.750 302.000 132.250 ;
        RECT 302.250 131.750 304.500 132.250 ;
        RECT 304.750 131.750 306.250 132.250 ;
        RECT 306.500 131.750 308.000 132.250 ;
        RECT 308.250 131.750 309.750 132.250 ;
        RECT 310.000 131.750 312.410 132.250 ;
        RECT 300.500 131.545 302.000 131.750 ;
        RECT 304.270 131.545 304.500 131.750 ;
        RECT 306.020 131.545 306.250 131.750 ;
        RECT 307.770 131.545 308.000 131.750 ;
        RECT 309.520 131.545 309.750 131.750 ;
        RECT 300.500 131.250 302.225 131.545 ;
        RECT 301.770 131.095 302.225 131.250 ;
        RECT 304.270 131.095 304.725 131.545 ;
        RECT 306.020 131.095 306.475 131.545 ;
        RECT 307.770 131.095 308.225 131.545 ;
        RECT 309.520 131.095 309.975 131.545 ;
        RECT 312.180 131.095 312.410 131.750 ;
        RECT 312.550 131.075 312.780 132.365 ;
        RECT 312.980 131.335 313.210 132.770 ;
        RECT 314.000 132.500 316.500 132.770 ;
        RECT 316.000 132.335 316.500 132.500 ;
        RECT 316.735 132.495 316.965 133.630 ;
        RECT 317.585 133.260 318.755 133.490 ;
        RECT 317.105 132.660 318.315 133.120 ;
        RECT 317.105 132.335 317.565 132.660 ;
        RECT 319.375 132.495 319.605 133.630 ;
        RECT 319.750 132.335 320.250 132.750 ;
        RECT 321.020 132.495 321.475 133.395 ;
        RECT 321.020 132.335 321.250 132.495 ;
        RECT 314.000 132.250 314.520 132.305 ;
        RECT 314.000 131.750 315.500 132.250 ;
        RECT 316.000 132.105 317.565 132.335 ;
        RECT 316.000 131.750 316.750 132.105 ;
        RECT 317.750 131.965 318.250 132.250 ;
        RECT 318.455 132.105 321.270 132.335 ;
        RECT 323.770 132.250 324.000 133.395 ;
        RECT 324.790 133.000 325.020 133.860 ;
        RECT 325.640 133.750 327.750 133.860 ;
        RECT 325.640 133.630 328.000 133.750 ;
        RECT 326.430 133.200 326.660 133.630 ;
        RECT 327.250 133.250 328.000 133.630 ;
        RECT 329.735 133.630 331.035 133.860 ;
        RECT 331.485 133.630 332.605 133.860 ;
        RECT 324.790 132.770 327.900 133.000 ;
        RECT 326.500 132.500 327.900 132.770 ;
        RECT 329.735 132.495 329.965 133.630 ;
        RECT 330.585 133.260 331.755 133.490 ;
        RECT 330.105 132.660 331.315 133.120 ;
        RECT 330.105 132.335 330.565 132.660 ;
        RECT 332.375 132.495 332.605 133.630 ;
        RECT 332.750 132.335 333.250 132.750 ;
        RECT 334.020 132.495 334.475 133.395 ;
        RECT 334.020 132.335 334.250 132.495 ;
        RECT 317.085 131.735 320.250 131.965 ;
        RECT 320.750 131.750 321.250 132.105 ;
        RECT 321.500 132.020 324.000 132.250 ;
        RECT 324.140 132.060 325.810 132.290 ;
        RECT 321.500 131.750 322.000 132.020 ;
        RECT 323.500 131.750 324.000 132.020 ;
        RECT 326.020 131.920 326.250 132.320 ;
        RECT 329.250 132.250 330.565 132.335 ;
        RECT 313.350 131.270 314.500 131.500 ;
        RECT 295.100 130.640 298.400 130.870 ;
        RECT 312.550 130.845 313.830 131.075 ;
        RECT 314.000 131.000 314.500 131.270 ;
        RECT 316.775 131.240 317.005 131.545 ;
        RECT 316.775 131.010 318.655 131.240 ;
        RECT 319.335 130.870 319.565 131.545 ;
        RECT 319.750 131.250 320.250 131.735 ;
        RECT 321.020 131.545 321.250 131.750 ;
        RECT 321.020 131.095 321.475 131.545 ;
        RECT 323.770 131.095 324.000 131.750 ;
        RECT 325.020 131.690 326.250 131.920 ;
        RECT 327.250 131.750 327.750 132.250 ;
        RECT 328.000 132.105 330.565 132.250 ;
        RECT 328.000 131.750 329.750 132.105 ;
        RECT 330.750 131.965 331.250 132.250 ;
        RECT 331.455 132.105 334.270 132.335 ;
        RECT 336.770 132.250 337.000 133.395 ;
        RECT 337.790 133.000 338.020 133.860 ;
        RECT 338.640 133.750 340.750 133.860 ;
        RECT 338.640 133.630 341.000 133.750 ;
        RECT 339.430 133.200 339.660 133.630 ;
        RECT 340.250 133.250 341.000 133.630 ;
        RECT 337.790 132.770 341.500 133.000 ;
        RECT 339.000 132.500 341.500 132.770 ;
        RECT 330.085 131.735 333.250 131.965 ;
        RECT 333.750 131.750 334.250 132.105 ;
        RECT 334.500 132.020 337.000 132.250 ;
        RECT 337.140 132.060 338.810 132.290 ;
        RECT 334.500 131.750 335.000 132.020 ;
        RECT 336.500 131.750 337.000 132.020 ;
        RECT 339.020 131.920 339.250 132.320 ;
        RECT 324.520 131.315 326.240 131.545 ;
        RECT 326.480 131.315 327.520 131.545 ;
        RECT 326.010 131.095 326.240 131.315 ;
        RECT 327.290 131.095 327.520 131.315 ;
        RECT 329.775 131.240 330.005 131.545 ;
        RECT 329.775 131.010 331.655 131.240 ;
        RECT 332.335 130.870 332.565 131.545 ;
        RECT 332.750 131.250 333.250 131.735 ;
        RECT 334.020 131.545 334.250 131.750 ;
        RECT 334.020 131.095 334.475 131.545 ;
        RECT 336.770 131.095 337.000 131.750 ;
        RECT 338.020 131.690 339.250 131.920 ;
        RECT 340.250 131.750 340.750 132.250 ;
        RECT 337.520 131.315 339.240 131.545 ;
        RECT 339.480 131.315 340.520 131.545 ;
        RECT 339.010 131.095 339.240 131.315 ;
        RECT 340.290 131.095 340.520 131.315 ;
        RECT 341.000 131.250 341.500 132.500 ;
        RECT 342.775 132.495 343.230 133.395 ;
        RECT 343.000 132.250 343.230 132.495 ;
        RECT 342.250 131.750 342.750 132.250 ;
        RECT 343.000 131.935 343.500 132.250 ;
        RECT 343.750 132.075 344.250 132.750 ;
        RECT 344.400 132.495 344.980 133.395 ;
        RECT 346.025 132.495 346.480 133.395 ;
        RECT 347.525 132.495 347.980 133.395 ;
        RECT 349.750 132.500 350.750 133.500 ;
        RECT 350.025 132.495 350.480 132.500 ;
        RECT 344.750 132.250 344.980 132.495 ;
        RECT 346.250 132.250 346.480 132.495 ;
        RECT 347.750 132.250 347.980 132.495 ;
        RECT 350.250 132.250 350.480 132.495 ;
        RECT 343.000 131.545 344.400 131.935 ;
        RECT 338.970 130.870 339.530 130.900 ;
        RECT 340.750 130.870 341.500 131.250 ;
        RECT 342.775 131.250 344.400 131.545 ;
        RECT 344.750 131.750 346.000 132.250 ;
        RECT 346.250 131.750 347.500 132.250 ;
        RECT 347.750 131.750 350.000 132.250 ;
        RECT 350.250 131.750 350.750 132.250 ;
        RECT 342.775 131.095 343.230 131.250 ;
        RECT 344.750 131.095 345.030 131.750 ;
        RECT 346.250 131.545 346.480 131.750 ;
        RECT 347.750 131.545 347.980 131.750 ;
        RECT 350.250 131.545 350.480 131.750 ;
        RECT 346.025 131.095 346.480 131.545 ;
        RECT 347.525 131.095 347.980 131.545 ;
        RECT 350.025 131.095 350.480 131.545 ;
        RECT 317.825 130.640 319.565 130.870 ;
        RECT 324.600 130.640 327.900 130.870 ;
        RECT 330.825 130.640 332.565 130.870 ;
        RECT 337.600 130.640 341.500 130.870 ;
        RECT 353.750 130.500 354.750 137.000 ;
        RECT 387.500 135.250 388.500 138.500 ;
        RECT 389.500 137.750 390.000 138.250 ;
        RECT 388.750 136.500 389.290 137.500 ;
        RECT 389.500 136.500 390.000 137.500 ;
        RECT 390.210 136.500 390.750 137.500 ;
        RECT 388.750 136.000 389.250 136.500 ;
        RECT 389.500 135.750 390.000 136.250 ;
        RECT 390.250 136.000 390.750 136.500 ;
        RECT 391.000 135.250 392.000 138.500 ;
        RECT 367.500 134.750 381.750 135.250 ;
        RECT 387.500 134.750 392.000 135.250 ;
        RECT 387.500 131.500 388.500 134.750 ;
        RECT 389.500 134.000 390.000 134.500 ;
        RECT 388.750 132.750 389.290 133.750 ;
        RECT 389.500 132.750 390.000 133.750 ;
        RECT 390.210 132.750 390.750 133.750 ;
        RECT 388.750 132.250 389.250 132.750 ;
        RECT 389.500 132.000 390.000 132.500 ;
        RECT 390.250 132.250 390.750 132.750 ;
        RECT 391.000 131.500 392.000 134.750 ;
        RECT 369.500 131.000 381.750 131.500 ;
        RECT 387.500 131.000 392.000 131.500 ;
        RECT 286.000 130.000 354.750 130.500 ;
        RECT 286.000 127.500 287.000 130.000 ;
        RECT 319.750 129.250 327.750 129.750 ;
        RECT 332.750 129.250 340.750 129.750 ;
        RECT 316.500 128.500 324.000 129.000 ;
        RECT 326.500 128.500 337.000 129.000 ;
        RECT 315.750 127.750 328.500 128.250 ;
        RECT 353.750 127.500 354.750 130.000 ;
        RECT 387.500 127.750 388.500 131.000 ;
        RECT 389.500 130.250 390.000 130.750 ;
        RECT 388.750 129.000 389.290 130.000 ;
        RECT 389.500 129.000 390.000 130.000 ;
        RECT 390.210 129.000 390.750 130.000 ;
        RECT 388.750 128.500 389.250 129.000 ;
        RECT 389.500 128.250 390.000 128.750 ;
        RECT 390.250 128.500 390.750 129.000 ;
        RECT 391.000 127.750 392.000 131.000 ;
        RECT 286.000 126.500 354.750 127.500 ;
        RECT 371.500 127.250 381.750 127.750 ;
        RECT 387.500 127.250 392.000 127.750 ;
        RECT 294.000 125.500 350.500 126.500 ;
        RECT 294.000 120.250 295.000 125.500 ;
        RECT 301.750 124.500 312.500 125.000 ;
        RECT 312.750 124.500 326.000 125.000 ;
        RECT 327.750 124.500 342.000 125.000 ;
        RECT 295.500 123.750 347.500 124.250 ;
        RECT 298.720 123.350 300.910 123.580 ;
        RECT 309.720 123.350 311.910 123.580 ;
        RECT 314.720 123.350 316.910 123.580 ;
        RECT 325.720 123.350 327.910 123.580 ;
        RECT 330.720 123.350 332.910 123.580 ;
        RECT 341.720 123.350 343.910 123.580 ;
        RECT 300.250 122.750 300.750 123.350 ;
        RECT 298.840 122.250 302.250 122.750 ;
        RECT 299.000 121.500 300.000 122.000 ;
        RECT 300.250 120.665 300.750 122.250 ;
        RECT 302.490 122.000 302.720 123.145 ;
        RECT 304.275 122.500 304.730 123.145 ;
        RECT 306.410 122.500 306.640 123.145 ;
        RECT 308.910 122.500 309.140 123.145 ;
        RECT 311.250 122.750 311.750 123.350 ;
        RECT 304.275 122.245 306.000 122.500 ;
        RECT 304.500 122.000 306.000 122.245 ;
        RECT 302.490 121.500 304.250 122.000 ;
        RECT 304.500 121.500 305.000 122.000 ;
        RECT 305.500 121.855 306.000 122.000 ;
        RECT 306.250 122.000 307.500 122.500 ;
        RECT 306.250 121.855 306.750 122.000 ;
        RECT 305.500 121.500 306.650 121.685 ;
        RECT 302.050 120.845 302.280 121.295 ;
        RECT 302.490 120.845 302.720 121.500 ;
        RECT 304.500 121.295 304.730 121.500 ;
        RECT 304.275 120.845 304.730 121.295 ;
        RECT 305.250 121.455 306.650 121.500 ;
        RECT 307.000 121.500 307.500 122.000 ;
        RECT 308.000 121.855 308.500 122.500 ;
        RECT 308.750 122.055 309.250 122.500 ;
        RECT 309.500 122.250 311.750 122.750 ;
        RECT 308.750 121.825 310.500 122.055 ;
        RECT 308.000 121.500 309.150 121.685 ;
        RECT 310.000 121.500 310.500 121.825 ;
        RECT 307.000 121.455 309.150 121.500 ;
        RECT 305.250 121.000 306.000 121.455 ;
        RECT 307.000 121.000 308.500 121.455 ;
        RECT 311.250 120.665 311.750 122.250 ;
        RECT 313.490 122.000 313.720 123.145 ;
        RECT 316.250 122.750 316.750 123.350 ;
        RECT 314.840 122.250 318.250 122.750 ;
        RECT 313.490 121.500 314.000 122.000 ;
        RECT 315.000 121.500 316.000 122.000 ;
        RECT 313.050 120.845 313.280 121.295 ;
        RECT 313.490 120.845 313.720 121.500 ;
        RECT 316.250 120.665 316.750 122.250 ;
        RECT 318.490 122.000 318.720 123.145 ;
        RECT 320.275 122.500 320.730 123.145 ;
        RECT 322.410 122.500 322.640 123.145 ;
        RECT 324.910 122.500 325.140 123.145 ;
        RECT 327.250 122.750 327.750 123.350 ;
        RECT 320.275 122.245 322.000 122.500 ;
        RECT 320.500 122.000 322.000 122.245 ;
        RECT 318.490 121.500 320.250 122.000 ;
        RECT 320.500 121.500 321.000 122.000 ;
        RECT 321.500 121.855 322.000 122.000 ;
        RECT 322.250 122.000 323.500 122.500 ;
        RECT 322.250 121.855 322.750 122.000 ;
        RECT 321.500 121.500 322.650 121.685 ;
        RECT 318.050 120.845 318.280 121.295 ;
        RECT 318.490 120.845 318.720 121.500 ;
        RECT 320.500 121.295 320.730 121.500 ;
        RECT 320.275 120.845 320.730 121.295 ;
        RECT 321.250 121.455 322.650 121.500 ;
        RECT 323.000 121.500 323.500 122.000 ;
        RECT 324.000 121.855 324.500 122.500 ;
        RECT 324.750 122.055 325.250 122.500 ;
        RECT 325.500 122.250 327.750 122.750 ;
        RECT 324.750 121.825 326.500 122.055 ;
        RECT 324.000 121.500 325.150 121.685 ;
        RECT 326.000 121.500 326.500 121.825 ;
        RECT 323.000 121.455 325.150 121.500 ;
        RECT 321.250 121.000 322.000 121.455 ;
        RECT 323.000 121.000 324.500 121.455 ;
        RECT 327.250 120.665 327.750 122.250 ;
        RECT 329.490 122.000 329.720 123.145 ;
        RECT 332.250 122.750 332.750 123.350 ;
        RECT 330.840 122.250 334.250 122.750 ;
        RECT 329.490 121.500 330.000 122.000 ;
        RECT 331.000 121.500 332.000 122.000 ;
        RECT 329.050 120.845 329.280 121.295 ;
        RECT 329.490 120.845 329.720 121.500 ;
        RECT 332.250 120.665 332.750 122.250 ;
        RECT 334.490 122.000 334.720 123.145 ;
        RECT 336.275 122.500 336.730 123.145 ;
        RECT 338.410 122.500 338.640 123.145 ;
        RECT 340.910 122.500 341.140 123.145 ;
        RECT 343.250 122.750 343.750 123.350 ;
        RECT 336.275 122.245 338.000 122.500 ;
        RECT 336.500 122.000 338.000 122.245 ;
        RECT 334.490 121.500 336.250 122.000 ;
        RECT 336.500 121.500 337.000 122.000 ;
        RECT 337.500 121.855 338.000 122.000 ;
        RECT 338.250 122.000 339.500 122.500 ;
        RECT 338.250 121.855 338.750 122.000 ;
        RECT 337.500 121.500 338.650 121.685 ;
        RECT 334.050 120.845 334.280 121.295 ;
        RECT 334.490 120.845 334.720 121.500 ;
        RECT 336.500 121.295 336.730 121.500 ;
        RECT 336.275 120.845 336.730 121.295 ;
        RECT 337.250 121.455 338.650 121.500 ;
        RECT 339.000 121.500 339.500 122.000 ;
        RECT 340.000 121.855 340.500 122.500 ;
        RECT 340.750 122.055 341.250 122.500 ;
        RECT 341.500 122.250 343.750 122.750 ;
        RECT 340.750 121.825 342.500 122.055 ;
        RECT 340.000 121.500 341.150 121.685 ;
        RECT 342.000 121.500 342.500 121.825 ;
        RECT 339.000 121.455 341.150 121.500 ;
        RECT 337.250 121.000 338.000 121.455 ;
        RECT 339.000 121.000 340.500 121.455 ;
        RECT 343.250 120.665 343.750 122.250 ;
        RECT 345.490 122.000 345.720 123.145 ;
        RECT 345.490 121.500 346.000 122.000 ;
        RECT 345.050 120.845 345.280 121.295 ;
        RECT 345.490 120.845 345.720 121.500 ;
        RECT 298.720 120.435 301.630 120.665 ;
        RECT 309.720 120.435 312.630 120.665 ;
        RECT 314.720 120.435 317.630 120.665 ;
        RECT 325.720 120.435 328.630 120.665 ;
        RECT 330.720 120.435 333.630 120.665 ;
        RECT 341.720 120.435 344.630 120.665 ;
        RECT 349.500 120.250 350.500 125.500 ;
        RECT 387.500 124.000 388.500 127.250 ;
        RECT 389.500 126.500 390.000 127.000 ;
        RECT 388.750 125.250 389.290 126.250 ;
        RECT 389.500 125.250 390.000 126.250 ;
        RECT 390.210 125.250 390.750 126.250 ;
        RECT 388.750 124.750 389.250 125.250 ;
        RECT 389.500 124.500 390.000 125.000 ;
        RECT 390.250 124.750 390.750 125.250 ;
        RECT 391.000 124.000 392.000 127.250 ;
        RECT 373.500 123.500 381.750 124.000 ;
        RECT 387.500 123.500 392.000 124.000 ;
        RECT 387.500 120.500 388.500 123.500 ;
        RECT 389.500 122.750 390.000 123.250 ;
        RECT 388.750 121.500 389.290 122.500 ;
        RECT 389.500 121.500 390.000 122.500 ;
        RECT 390.210 121.500 390.750 122.500 ;
        RECT 388.750 121.000 389.250 121.500 ;
        RECT 389.500 120.750 390.000 121.250 ;
        RECT 390.250 121.000 390.750 121.500 ;
        RECT 391.000 120.500 392.000 123.500 ;
        RECT 397.000 149.750 401.500 150.500 ;
        RECT 397.000 146.500 398.000 149.750 ;
        RECT 399.000 149.000 399.500 149.500 ;
        RECT 398.250 147.750 398.790 148.750 ;
        RECT 399.000 147.750 399.500 148.750 ;
        RECT 399.710 147.750 400.250 148.750 ;
        RECT 398.250 147.250 398.750 147.750 ;
        RECT 399.000 147.000 399.500 147.500 ;
        RECT 399.750 147.250 400.250 147.750 ;
        RECT 400.500 146.500 401.500 149.750 ;
        RECT 397.000 146.000 401.500 146.500 ;
        RECT 397.000 142.750 398.000 146.000 ;
        RECT 399.000 145.250 399.500 145.750 ;
        RECT 398.250 144.000 398.790 145.000 ;
        RECT 399.000 144.000 399.500 145.000 ;
        RECT 399.710 144.000 400.250 145.000 ;
        RECT 398.250 143.500 398.750 144.000 ;
        RECT 399.000 143.250 399.500 143.750 ;
        RECT 399.750 143.500 400.250 144.000 ;
        RECT 400.500 142.750 401.500 146.000 ;
        RECT 397.000 142.250 401.500 142.750 ;
        RECT 397.000 139.000 398.000 142.250 ;
        RECT 399.000 141.500 399.500 142.000 ;
        RECT 398.250 140.250 398.790 141.250 ;
        RECT 399.000 140.250 399.500 141.250 ;
        RECT 399.710 140.250 400.250 141.250 ;
        RECT 398.250 139.750 398.750 140.250 ;
        RECT 399.000 139.500 399.500 140.000 ;
        RECT 399.750 139.750 400.250 140.250 ;
        RECT 400.500 139.000 401.500 142.250 ;
        RECT 397.000 138.500 401.500 139.000 ;
        RECT 397.000 135.250 398.000 138.500 ;
        RECT 399.000 137.750 399.500 138.250 ;
        RECT 398.250 136.500 398.790 137.500 ;
        RECT 399.000 136.500 399.500 137.500 ;
        RECT 399.710 136.500 400.250 137.500 ;
        RECT 398.250 136.000 398.750 136.500 ;
        RECT 399.000 135.750 399.500 136.250 ;
        RECT 399.750 136.000 400.250 136.500 ;
        RECT 400.500 135.250 401.500 138.500 ;
        RECT 397.000 134.750 401.500 135.250 ;
        RECT 397.000 131.500 398.000 134.750 ;
        RECT 399.000 134.000 399.500 134.500 ;
        RECT 398.250 132.750 398.790 133.750 ;
        RECT 399.000 132.750 399.500 133.750 ;
        RECT 399.710 132.750 400.250 133.750 ;
        RECT 398.250 132.250 398.750 132.750 ;
        RECT 399.000 132.000 399.500 132.500 ;
        RECT 399.750 132.250 400.250 132.750 ;
        RECT 400.500 131.500 401.500 134.750 ;
        RECT 397.000 131.000 401.500 131.500 ;
        RECT 397.000 127.750 398.000 131.000 ;
        RECT 399.000 130.250 399.500 130.750 ;
        RECT 398.250 129.000 398.790 130.000 ;
        RECT 399.000 129.000 399.500 130.000 ;
        RECT 399.710 129.000 400.250 130.000 ;
        RECT 398.250 128.500 398.750 129.000 ;
        RECT 399.000 128.250 399.500 128.750 ;
        RECT 399.750 128.500 400.250 129.000 ;
        RECT 400.500 127.750 401.500 131.000 ;
        RECT 397.000 127.250 401.500 127.750 ;
        RECT 397.000 124.000 398.000 127.250 ;
        RECT 399.000 126.500 399.500 127.000 ;
        RECT 398.250 125.250 398.790 126.250 ;
        RECT 399.000 125.250 399.500 126.250 ;
        RECT 399.710 125.250 400.250 126.250 ;
        RECT 398.250 124.750 398.750 125.250 ;
        RECT 399.000 124.500 399.500 125.000 ;
        RECT 399.750 124.750 400.250 125.250 ;
        RECT 400.500 124.000 401.500 127.250 ;
        RECT 397.000 123.500 401.500 124.000 ;
        RECT 397.000 120.500 398.000 123.500 ;
        RECT 399.000 122.750 399.500 123.250 ;
        RECT 398.250 121.500 398.790 122.500 ;
        RECT 399.000 121.500 399.500 122.500 ;
        RECT 399.710 121.500 400.250 122.500 ;
        RECT 398.250 121.000 398.750 121.500 ;
        RECT 399.000 120.750 399.500 121.250 ;
        RECT 399.750 121.000 400.250 121.500 ;
        RECT 400.500 120.500 401.500 123.500 ;
        RECT 406.500 149.750 411.000 150.500 ;
        RECT 406.500 146.500 407.500 149.750 ;
        RECT 408.500 149.000 409.000 149.500 ;
        RECT 407.750 147.750 408.290 148.750 ;
        RECT 408.500 147.750 409.000 148.750 ;
        RECT 409.210 147.750 409.750 148.750 ;
        RECT 407.750 147.250 408.250 147.750 ;
        RECT 408.500 147.000 409.000 147.500 ;
        RECT 409.250 147.250 409.750 147.750 ;
        RECT 410.000 146.500 411.000 149.750 ;
        RECT 406.500 146.000 411.000 146.500 ;
        RECT 406.500 142.750 407.500 146.000 ;
        RECT 408.500 145.250 409.000 145.750 ;
        RECT 407.750 144.000 408.290 145.000 ;
        RECT 408.500 144.000 409.000 145.000 ;
        RECT 409.210 144.000 409.750 145.000 ;
        RECT 407.750 143.500 408.250 144.000 ;
        RECT 408.500 143.250 409.000 143.750 ;
        RECT 409.250 143.500 409.750 144.000 ;
        RECT 410.000 142.750 411.000 146.000 ;
        RECT 406.500 142.250 411.000 142.750 ;
        RECT 406.500 139.000 407.500 142.250 ;
        RECT 408.500 141.500 409.000 142.000 ;
        RECT 407.750 140.250 408.290 141.250 ;
        RECT 408.500 140.250 409.000 141.250 ;
        RECT 409.210 140.250 409.750 141.250 ;
        RECT 407.750 139.750 408.250 140.250 ;
        RECT 408.500 139.500 409.000 140.000 ;
        RECT 409.250 139.750 409.750 140.250 ;
        RECT 410.000 139.000 411.000 142.250 ;
        RECT 406.500 138.500 411.000 139.000 ;
        RECT 406.500 135.250 407.500 138.500 ;
        RECT 408.500 137.750 409.000 138.250 ;
        RECT 407.750 136.500 408.290 137.500 ;
        RECT 408.500 136.500 409.000 137.500 ;
        RECT 409.210 136.500 409.750 137.500 ;
        RECT 407.750 136.000 408.250 136.500 ;
        RECT 408.500 135.750 409.000 136.250 ;
        RECT 409.250 136.000 409.750 136.500 ;
        RECT 410.000 135.250 411.000 138.500 ;
        RECT 406.500 134.750 411.000 135.250 ;
        RECT 406.500 131.500 407.500 134.750 ;
        RECT 408.500 134.000 409.000 134.500 ;
        RECT 407.750 132.750 408.290 133.750 ;
        RECT 408.500 132.750 409.000 133.750 ;
        RECT 409.210 132.750 409.750 133.750 ;
        RECT 407.750 132.250 408.250 132.750 ;
        RECT 408.500 132.000 409.000 132.500 ;
        RECT 409.250 132.250 409.750 132.750 ;
        RECT 410.000 131.500 411.000 134.750 ;
        RECT 406.500 131.000 411.000 131.500 ;
        RECT 406.500 127.750 407.500 131.000 ;
        RECT 408.500 130.250 409.000 130.750 ;
        RECT 407.750 129.000 408.290 130.000 ;
        RECT 408.500 129.000 409.000 130.000 ;
        RECT 409.210 129.000 409.750 130.000 ;
        RECT 407.750 128.500 408.250 129.000 ;
        RECT 408.500 128.250 409.000 128.750 ;
        RECT 409.250 128.500 409.750 129.000 ;
        RECT 410.000 127.750 411.000 131.000 ;
        RECT 406.500 127.250 411.000 127.750 ;
        RECT 406.500 124.000 407.500 127.250 ;
        RECT 408.500 126.500 409.000 127.000 ;
        RECT 407.750 125.250 408.290 126.250 ;
        RECT 408.500 125.250 409.000 126.250 ;
        RECT 409.210 125.250 409.750 126.250 ;
        RECT 407.750 124.750 408.250 125.250 ;
        RECT 408.500 124.500 409.000 125.000 ;
        RECT 409.250 124.750 409.750 125.250 ;
        RECT 410.000 124.000 411.000 127.250 ;
        RECT 406.500 123.500 411.000 124.000 ;
        RECT 406.500 120.500 407.500 123.500 ;
        RECT 408.500 122.750 409.000 123.250 ;
        RECT 407.750 121.500 408.290 122.500 ;
        RECT 408.500 121.500 409.000 122.500 ;
        RECT 409.210 121.500 409.750 122.500 ;
        RECT 407.750 121.000 408.250 121.500 ;
        RECT 408.500 120.750 409.000 121.250 ;
        RECT 409.250 121.000 409.750 121.500 ;
        RECT 410.000 120.500 411.000 123.500 ;
        RECT 294.000 119.750 350.500 120.250 ;
        RECT 294.000 114.000 295.000 119.750 ;
        RECT 299.500 119.000 314.000 119.500 ;
        RECT 315.500 119.000 330.000 119.500 ;
        RECT 331.500 119.000 346.000 119.500 ;
        RECT 298.750 118.250 313.250 118.750 ;
        RECT 314.750 118.250 321.750 118.750 ;
        RECT 322.000 118.250 330.500 118.750 ;
        RECT 330.750 118.250 337.750 118.750 ;
        RECT 338.000 118.250 344.000 118.750 ;
        RECT 295.500 117.500 347.500 118.000 ;
        RECT 301.220 117.100 303.410 117.330 ;
        RECT 308.220 117.100 310.410 117.330 ;
        RECT 317.220 117.100 319.410 117.330 ;
        RECT 321.970 117.100 324.160 117.330 ;
        RECT 333.220 117.100 335.410 117.330 ;
        RECT 339.720 117.100 341.910 117.330 ;
        RECT 299.275 115.995 299.730 116.895 ;
        RECT 301.340 116.000 302.000 116.500 ;
        RECT 299.500 115.750 299.730 115.995 ;
        RECT 304.990 115.750 305.220 116.895 ;
        RECT 307.250 116.500 308.250 116.750 ;
        RECT 307.250 116.000 309.500 116.500 ;
        RECT 307.250 115.750 308.250 116.000 ;
        RECT 311.990 115.750 312.220 116.895 ;
        RECT 315.275 115.995 315.730 116.895 ;
        RECT 320.990 116.500 321.220 116.895 ;
        RECT 317.340 116.000 318.000 116.500 ;
        RECT 320.990 116.000 322.750 116.500 ;
        RECT 315.500 115.750 315.730 115.995 ;
        RECT 298.750 115.250 299.250 115.750 ;
        RECT 299.500 115.250 302.000 115.750 ;
        RECT 304.990 115.250 305.750 115.750 ;
        RECT 308.560 115.405 311.850 115.635 ;
        RECT 311.990 115.250 312.500 115.750 ;
        RECT 314.750 115.250 315.250 115.750 ;
        RECT 315.500 115.250 318.000 115.750 ;
        RECT 320.990 115.250 321.750 116.000 ;
        RECT 325.740 115.750 325.970 116.895 ;
        RECT 328.275 115.995 328.730 116.895 ;
        RECT 329.775 115.995 330.230 116.895 ;
        RECT 331.275 115.995 331.730 116.895 ;
        RECT 336.990 116.500 337.220 116.895 ;
        RECT 333.340 116.000 334.000 116.500 ;
        RECT 336.990 116.000 340.500 116.500 ;
        RECT 328.500 115.750 328.730 115.995 ;
        RECT 330.000 115.750 330.230 115.995 ;
        RECT 331.500 115.750 331.730 115.995 ;
        RECT 322.310 115.405 325.600 115.635 ;
        RECT 325.740 115.250 328.250 115.750 ;
        RECT 328.500 115.250 329.750 115.750 ;
        RECT 330.000 115.250 330.500 115.750 ;
        RECT 330.750 115.250 331.250 115.750 ;
        RECT 331.500 115.250 334.000 115.750 ;
        RECT 336.990 115.250 337.750 116.000 ;
        RECT 343.490 115.750 343.720 116.895 ;
        RECT 340.060 115.405 343.350 115.635 ;
        RECT 343.490 115.250 344.000 115.750 ;
        RECT 299.500 115.045 299.730 115.250 ;
        RECT 299.275 114.595 299.730 115.045 ;
        RECT 304.550 114.595 304.780 115.045 ;
        RECT 304.990 114.595 305.220 115.250 ;
        RECT 311.550 114.595 311.780 115.045 ;
        RECT 311.990 114.595 312.220 115.250 ;
        RECT 315.500 115.045 315.730 115.250 ;
        RECT 315.275 114.595 315.730 115.045 ;
        RECT 320.550 114.595 320.780 115.045 ;
        RECT 320.990 114.595 321.220 115.250 ;
        RECT 325.300 114.595 325.530 115.045 ;
        RECT 325.740 114.595 325.970 115.250 ;
        RECT 328.500 115.045 328.730 115.250 ;
        RECT 330.000 115.045 330.230 115.250 ;
        RECT 331.500 115.045 331.730 115.250 ;
        RECT 328.275 114.595 328.730 115.045 ;
        RECT 329.775 114.595 330.230 115.045 ;
        RECT 331.275 114.595 331.730 115.045 ;
        RECT 336.550 114.595 336.780 115.045 ;
        RECT 336.990 114.595 337.220 115.250 ;
        RECT 343.050 114.595 343.280 115.045 ;
        RECT 343.490 114.595 343.720 115.250 ;
        RECT 301.220 114.185 304.130 114.415 ;
        RECT 308.220 114.185 311.130 114.415 ;
        RECT 317.220 114.185 320.130 114.415 ;
        RECT 321.970 114.185 324.880 114.415 ;
        RECT 333.220 114.185 336.130 114.415 ;
        RECT 339.720 114.185 342.630 114.415 ;
        RECT 349.500 114.000 350.500 119.750 ;
        RECT 382.750 119.500 411.250 120.500 ;
        RECT 294.000 113.500 350.500 114.000 ;
        RECT 294.000 113.000 295.000 113.500 ;
        RECT 349.500 113.000 350.500 113.500 ;
        RECT 284.500 109.000 425.000 113.000 ;
        RECT 284.500 104.000 425.000 108.000 ;
      LAYER met2 ;
        RECT 285.500 104.000 286.750 204.000 ;
        RECT 287.750 109.000 289.000 209.000 ;
        RECT 290.000 158.500 291.000 204.000 ;
        RECT 291.500 158.500 292.500 209.000 ;
        RECT 296.790 182.765 297.070 183.135 ;
        RECT 300.485 182.765 300.765 183.135 ;
        RECT 296.330 181.265 296.610 181.635 ;
        RECT 296.400 176.550 296.540 181.265 ;
        RECT 296.860 176.890 297.000 182.765 ;
        RECT 297.710 181.265 297.990 181.635 ;
        RECT 297.260 179.290 297.520 179.610 ;
        RECT 297.320 178.635 297.460 179.290 ;
        RECT 297.250 178.265 297.530 178.635 ;
        RECT 296.800 176.570 297.060 176.890 ;
        RECT 296.340 176.230 296.600 176.550 ;
        RECT 295.880 175.890 296.140 176.210 ;
        RECT 295.420 170.110 295.680 170.430 ;
        RECT 295.480 165.135 295.620 170.110 ;
        RECT 295.940 168.135 296.080 175.890 ;
        RECT 296.400 173.830 296.540 176.230 ;
        RECT 296.860 176.210 297.000 176.570 ;
        RECT 296.800 175.890 297.060 176.210 ;
        RECT 296.340 173.510 296.600 173.830 ;
        RECT 296.400 170.770 296.540 173.510 ;
        RECT 296.860 171.790 297.000 175.890 ;
        RECT 297.320 175.870 297.460 178.265 ;
        RECT 297.780 176.550 297.920 181.265 ;
        RECT 300.010 179.765 300.290 180.135 ;
        RECT 299.100 179.290 299.360 179.610 ;
        RECT 300.080 179.270 300.220 179.765 ;
        RECT 300.020 178.950 300.280 179.270 ;
        RECT 298.180 178.270 298.440 178.590 ;
        RECT 297.720 176.230 297.980 176.550 ;
        RECT 297.260 175.550 297.520 175.870 ;
        RECT 297.320 174.170 297.460 175.550 ;
        RECT 297.260 173.850 297.520 174.170 ;
        RECT 297.780 173.150 297.920 176.230 ;
        RECT 298.240 176.210 298.380 178.270 ;
        RECT 300.080 177.230 300.220 178.950 ;
        RECT 300.555 177.570 300.695 182.765 ;
        RECT 311.870 180.455 313.410 180.825 ;
        RECT 300.960 179.765 301.240 180.135 ;
        RECT 312.440 179.970 312.700 180.290 ;
        RECT 312.900 179.970 313.160 180.290 ;
        RECT 300.495 177.250 300.755 177.570 ;
        RECT 300.020 176.910 300.280 177.230 ;
        RECT 298.180 175.890 298.440 176.210 ;
        RECT 297.720 172.830 297.980 173.150 ;
        RECT 296.800 171.470 297.060 171.790 ;
        RECT 296.340 170.450 296.600 170.770 ;
        RECT 295.870 167.765 296.150 168.135 ;
        RECT 295.410 164.765 295.690 165.135 ;
        RECT 296.860 163.630 297.000 171.470 ;
        RECT 298.240 171.450 298.380 175.890 ;
        RECT 299.560 173.850 299.820 174.170 ;
        RECT 298.640 173.170 298.900 173.490 ;
        RECT 297.720 171.130 297.980 171.450 ;
        RECT 298.180 171.130 298.440 171.450 ;
        RECT 297.780 166.635 297.920 171.130 ;
        RECT 298.180 170.450 298.440 170.770 ;
        RECT 297.710 166.265 297.990 166.635 ;
        RECT 297.260 165.690 297.520 166.010 ;
        RECT 296.800 163.310 297.060 163.630 ;
        RECT 297.320 163.290 297.460 165.690 ;
        RECT 298.240 164.990 298.380 170.450 ;
        RECT 298.700 166.690 298.840 173.170 ;
        RECT 298.640 166.370 298.900 166.690 ;
        RECT 298.700 165.330 298.840 166.370 ;
        RECT 299.620 165.330 299.760 173.850 ;
        RECT 300.080 173.490 300.220 176.910 ;
        RECT 300.020 173.170 300.280 173.490 ;
        RECT 300.480 165.350 300.740 165.670 ;
        RECT 298.640 165.010 298.900 165.330 ;
        RECT 299.560 165.010 299.820 165.330 ;
        RECT 298.180 164.670 298.440 164.990 ;
        RECT 298.240 163.970 298.380 164.670 ;
        RECT 298.180 163.650 298.440 163.970 ;
        RECT 300.540 163.735 300.680 165.350 ;
        RECT 300.470 163.365 300.750 163.735 ;
        RECT 297.260 162.970 297.520 163.290 ;
        RECT 300.480 162.970 300.740 163.365 ;
        RECT 299.560 162.290 299.820 162.610 ;
        RECT 294.500 161.950 294.760 162.270 ;
        RECT 296.340 161.950 296.600 162.270 ;
        RECT 299.620 162.135 299.760 162.290 ;
        RECT 301.030 162.270 301.170 179.765 ;
        RECT 310.600 179.630 310.860 179.950 ;
        RECT 301.435 178.265 301.715 178.635 ;
        RECT 301.505 166.010 301.645 178.265 ;
        RECT 310.660 170.770 310.800 179.630 ;
        RECT 311.060 179.290 311.320 179.610 ;
        RECT 311.120 177.230 311.260 179.290 ;
        RECT 311.060 176.910 311.320 177.230 ;
        RECT 311.120 171.110 311.260 176.910 ;
        RECT 312.500 176.210 312.640 179.970 ;
        RECT 312.960 177.570 313.100 179.970 ;
        RECT 314.740 178.610 315.000 178.930 ;
        RECT 312.900 177.250 313.160 177.570 ;
        RECT 313.810 176.765 314.090 177.135 ;
        RECT 312.440 175.890 312.700 176.210 ;
        RECT 312.900 175.550 313.160 175.870 ;
        RECT 312.960 171.110 313.100 175.550 ;
        RECT 313.350 172.265 313.630 172.635 ;
        RECT 311.060 170.790 311.320 171.110 ;
        RECT 312.900 170.790 313.160 171.110 ;
        RECT 310.600 170.450 310.860 170.770 ;
        RECT 301.445 165.690 301.705 166.010 ;
        RECT 310.660 163.290 310.800 170.450 ;
        RECT 311.120 168.730 311.260 170.790 ;
        RECT 312.960 169.635 313.100 170.790 ;
        RECT 312.890 169.265 313.170 169.635 ;
        RECT 311.060 168.410 311.320 168.730 ;
        RECT 313.420 168.050 313.560 172.265 ;
        RECT 313.360 167.730 313.620 168.050 ;
        RECT 311.520 165.010 311.780 165.330 ;
        RECT 311.580 163.970 311.720 165.010 ;
        RECT 311.520 163.650 311.780 163.970 ;
        RECT 310.600 162.970 310.860 163.290 ;
        RECT 313.880 162.610 314.020 176.765 ;
        RECT 314.270 175.265 314.550 175.635 ;
        RECT 314.340 166.690 314.480 175.265 ;
        RECT 314.800 174.135 314.940 178.610 ;
        RECT 314.730 173.765 315.010 174.135 ;
        RECT 317.030 170.765 317.310 171.135 ;
        RECT 317.040 170.450 317.300 170.765 ;
        RECT 314.280 166.370 314.540 166.690 ;
        RECT 314.340 163.290 314.480 166.370 ;
        RECT 314.280 162.970 314.540 163.290 ;
        RECT 313.820 162.290 314.080 162.610 ;
        RECT 294.560 160.635 294.700 161.950 ;
        RECT 299.550 161.765 299.830 162.135 ;
        RECT 300.970 161.950 301.230 162.270 ;
        RECT 294.490 160.265 294.770 160.635 ;
        RECT 318.000 158.500 319.000 204.000 ;
        RECT 319.500 158.500 320.500 209.000 ;
        RECT 321.250 183.500 322.500 209.000 ;
        RECT 322.750 183.500 324.000 204.000 ;
        RECT 324.250 183.500 325.500 199.000 ;
        RECT 326.520 187.250 327.020 194.500 ;
        RECT 327.270 188.000 327.770 193.750 ;
        RECT 328.020 191.750 328.520 197.500 ;
        RECT 328.020 185.000 328.520 190.000 ;
        RECT 329.680 188.000 330.180 193.750 ;
        RECT 330.430 187.250 330.930 194.500 ;
        RECT 331.340 191.750 331.840 194.500 ;
        RECT 331.340 185.000 331.840 190.750 ;
        RECT 332.090 188.000 332.590 193.750 ;
        RECT 332.840 187.250 333.340 191.500 ;
        RECT 333.750 187.250 334.250 194.500 ;
        RECT 334.500 188.000 335.000 193.750 ;
        RECT 335.250 187.250 335.750 194.500 ;
        RECT 336.160 191.000 336.660 194.500 ;
        RECT 336.910 188.000 337.410 193.750 ;
        RECT 337.660 191.750 338.160 197.500 ;
        RECT 337.660 187.250 338.160 190.000 ;
        RECT 338.570 187.250 339.070 194.500 ;
        RECT 339.320 188.000 339.820 193.750 ;
        RECT 340.980 191.750 341.480 194.500 ;
        RECT 340.980 187.250 341.480 190.750 ;
        RECT 341.730 188.000 342.230 193.750 ;
        RECT 289.500 146.500 290.750 150.750 ;
        RECT 291.000 126.500 292.000 153.000 ;
        RECT 292.250 126.500 293.250 155.500 ;
        RECT 299.250 149.500 301.250 158.000 ;
        RECT 296.000 146.500 296.500 149.250 ;
        RECT 293.750 143.250 294.250 146.250 ;
        RECT 294.000 138.750 294.500 143.000 ;
        RECT 299.750 142.500 300.250 145.750 ;
        RECT 302.250 143.250 302.750 146.750 ;
        RECT 303.750 146.500 304.250 149.250 ;
        RECT 294.000 131.750 294.500 136.750 ;
        RECT 295.000 136.250 295.500 139.250 ;
        RECT 295.750 132.500 296.250 139.250 ;
        RECT 297.000 133.250 297.500 135.250 ;
        RECT 297.750 131.750 298.250 136.000 ;
        RECT 298.500 131.750 299.000 139.750 ;
        RECT 303.500 138.750 304.000 139.250 ;
        RECT 304.500 137.000 305.000 137.500 ;
        RECT 303.500 131.750 304.000 132.250 ;
        RECT 304.500 130.000 305.000 130.500 ;
        RECT 305.500 130.000 306.000 144.500 ;
        RECT 306.250 134.000 306.750 148.500 ;
        RECT 307.750 143.250 308.250 150.750 ;
        RECT 310.750 146.500 311.250 149.250 ;
        RECT 310.000 143.250 310.500 146.250 ;
        RECT 307.500 135.500 308.000 139.250 ;
        RECT 311.500 138.750 312.000 150.000 ;
        RECT 311.000 137.000 311.500 137.500 ;
        RECT 308.750 131.750 309.250 135.250 ;
        RECT 311.750 131.750 312.250 132.250 ;
        RECT 312.500 130.000 313.000 144.500 ;
        RECT 313.250 134.000 313.750 148.500 ;
        RECT 314.750 143.250 315.250 146.750 ;
        RECT 319.000 146.500 319.500 149.250 ;
        RECT 323.000 143.250 323.500 146.250 ;
        RECT 314.000 131.000 314.500 143.000 ;
        RECT 314.750 136.250 315.250 142.250 ;
        RECT 315.500 140.250 316.000 142.250 ;
        RECT 315.750 136.250 316.250 139.250 ;
        RECT 315.000 131.750 315.500 135.250 ;
        RECT 315.750 127.750 316.250 133.750 ;
        RECT 316.500 128.500 317.000 140.000 ;
        RECT 319.500 135.500 320.000 139.250 ;
        RECT 321.500 135.500 322.000 139.250 ;
        RECT 322.250 136.250 322.750 139.250 ;
        RECT 323.250 136.250 323.750 139.750 ;
        RECT 325.250 138.750 325.750 139.250 ;
        RECT 326.750 134.750 327.250 139.250 ;
        RECT 327.500 133.250 328.000 142.250 ;
        RECT 328.500 140.250 329.000 142.250 ;
        RECT 328.750 136.250 329.250 139.250 ;
        RECT 329.500 135.500 330.000 140.000 ;
        RECT 332.500 135.500 333.000 139.250 ;
        RECT 334.500 135.500 335.000 139.250 ;
        RECT 335.250 136.250 335.750 139.250 ;
        RECT 336.250 136.250 336.750 139.750 ;
        RECT 338.250 138.750 338.750 139.250 ;
        RECT 317.750 131.750 318.250 132.250 ;
        RECT 319.750 129.250 320.250 132.750 ;
        RECT 320.750 129.250 321.250 132.250 ;
        RECT 321.500 128.500 322.000 132.250 ;
        RECT 323.500 128.500 324.000 132.250 ;
        RECT 326.500 128.500 327.000 133.000 ;
        RECT 327.250 129.250 327.750 132.250 ;
        RECT 328.000 127.750 328.500 132.250 ;
        RECT 330.750 131.750 331.250 132.250 ;
        RECT 332.750 129.250 333.250 132.750 ;
        RECT 333.750 129.250 334.250 132.250 ;
        RECT 334.500 128.500 335.000 132.250 ;
        RECT 336.500 128.500 337.000 132.250 ;
        RECT 339.000 130.610 339.500 150.750 ;
        RECT 339.750 146.500 340.250 150.000 ;
        RECT 344.000 145.000 345.250 199.000 ;
        RECT 345.500 183.500 346.750 209.000 ;
        RECT 347.000 183.500 348.250 204.000 ;
        RECT 349.250 192.750 350.500 209.000 ;
        RECT 354.500 192.750 355.750 209.000 ;
        RECT 350.000 190.750 350.500 191.750 ;
        RECT 350.750 188.750 351.250 192.500 ;
        RECT 351.500 190.750 352.000 191.750 ;
        RECT 353.000 190.750 353.500 191.750 ;
        RECT 353.750 188.750 354.250 192.500 ;
        RECT 354.500 190.750 355.000 191.750 ;
        RECT 350.500 182.500 351.500 188.750 ;
        RECT 348.250 181.500 351.500 182.500 ;
        RECT 344.000 143.750 344.500 145.000 ;
        RECT 342.250 143.250 344.500 143.750 ;
        RECT 339.750 138.750 340.250 143.000 ;
        RECT 340.500 133.250 341.000 135.250 ;
        RECT 340.250 129.250 340.750 132.250 ;
        RECT 342.250 131.750 342.750 143.250 ;
        RECT 348.250 139.500 349.250 181.500 ;
        RECT 353.500 180.500 354.500 188.750 ;
        RECT 349.750 179.500 354.500 180.500 ;
        RECT 344.000 136.250 344.500 138.750 ;
        RECT 343.750 132.250 344.250 135.250 ;
        RECT 347.750 134.750 348.250 139.250 ;
        RECT 348.500 131.750 349.000 136.750 ;
        RECT 349.750 132.500 350.750 179.500 ;
        RECT 292.250 125.500 296.500 126.500 ;
        RECT 295.500 104.000 296.500 125.500 ;
        RECT 297.000 109.000 298.000 126.500 ;
        RECT 301.750 122.250 302.250 125.000 ;
        RECT 299.500 119.000 300.000 122.000 ;
        RECT 298.750 115.250 299.250 118.750 ;
        RECT 301.500 116.000 302.000 119.500 ;
        RECT 305.250 115.250 305.750 121.500 ;
        RECT 308.000 119.000 308.500 122.500 ;
        RECT 309.500 122.250 310.000 125.000 ;
        RECT 307.250 115.750 308.250 116.750 ;
        RECT 312.000 115.250 312.500 125.000 ;
        RECT 312.750 118.250 313.250 125.000 ;
        RECT 317.750 122.250 318.250 125.000 ;
        RECT 313.500 119.000 314.000 122.000 ;
        RECT 315.500 119.000 316.000 122.000 ;
        RECT 314.750 115.250 315.250 118.750 ;
        RECT 317.500 116.000 318.000 119.500 ;
        RECT 321.250 115.250 321.750 121.500 ;
        RECT 324.000 119.000 324.500 122.500 ;
        RECT 325.500 122.250 326.000 125.000 ;
        RECT 327.750 115.250 328.250 125.000 ;
        RECT 333.750 122.250 334.250 125.000 ;
        RECT 329.500 119.000 330.000 122.000 ;
        RECT 331.500 119.000 332.000 122.000 ;
        RECT 330.000 115.250 330.500 118.750 ;
        RECT 330.750 115.250 331.250 118.750 ;
        RECT 333.500 116.000 334.000 119.500 ;
        RECT 337.250 115.250 337.750 121.500 ;
        RECT 340.000 119.000 340.500 122.500 ;
        RECT 341.500 122.250 342.000 125.000 ;
        RECT 343.500 115.250 344.000 120.750 ;
        RECT 345.500 119.000 346.000 122.000 ;
        RECT 346.500 104.000 347.500 126.500 ;
        RECT 348.000 109.000 349.000 126.500 ;
        RECT 351.250 109.000 352.250 153.000 ;
        RECT 352.500 104.000 353.500 155.500 ;
        RECT 359.500 149.750 360.000 183.500 ;
        RECT 360.500 166.250 361.000 182.000 ;
        RECT 361.500 146.000 362.000 180.500 ;
        RECT 362.500 170.000 363.000 179.000 ;
        RECT 363.500 142.250 364.000 177.500 ;
        RECT 364.500 173.750 365.000 176.000 ;
        RECT 365.500 138.500 366.000 174.500 ;
        RECT 366.500 172.000 367.000 178.000 ;
        RECT 367.500 134.750 368.000 171.500 ;
        RECT 368.500 169.000 369.000 181.750 ;
        RECT 369.500 131.000 370.000 168.500 ;
        RECT 370.500 166.000 371.000 185.500 ;
        RECT 371.500 127.250 372.000 165.500 ;
        RECT 372.500 163.000 373.000 189.250 ;
        RECT 373.500 123.500 374.000 162.500 ;
        RECT 374.500 160.000 375.000 193.000 ;
        RECT 379.000 165.000 380.000 204.000 ;
        RECT 382.750 196.000 383.750 209.000 ;
        RECT 387.500 196.000 388.500 209.000 ;
        RECT 391.000 196.000 392.000 209.000 ;
        RECT 392.750 196.000 393.250 197.000 ;
        RECT 397.000 196.000 398.000 209.000 ;
        RECT 400.500 196.000 401.500 209.000 ;
        RECT 402.250 196.000 402.750 197.000 ;
        RECT 406.500 196.000 407.500 209.000 ;
        RECT 410.000 196.000 411.000 209.000 ;
        RECT 423.000 205.000 427.000 209.000 ;
        RECT 388.750 195.000 389.250 195.500 ;
        RECT 390.250 195.000 390.750 195.500 ;
        RECT 398.250 195.000 398.750 195.500 ;
        RECT 399.750 195.000 400.250 195.500 ;
        RECT 407.750 195.000 408.250 195.500 ;
        RECT 409.250 195.000 409.750 195.500 ;
        RECT 389.500 194.000 390.000 194.500 ;
        RECT 399.000 194.000 399.500 194.500 ;
        RECT 408.500 194.000 409.000 194.500 ;
        RECT 389.500 193.000 390.000 193.750 ;
        RECT 399.000 193.000 399.500 193.750 ;
        RECT 408.500 193.000 409.000 193.750 ;
        RECT 381.250 192.500 411.250 193.000 ;
        RECT 388.750 191.250 389.250 191.750 ;
        RECT 390.250 191.250 390.750 191.750 ;
        RECT 398.250 191.250 398.750 191.750 ;
        RECT 399.750 191.250 400.250 191.750 ;
        RECT 407.750 191.250 408.250 191.750 ;
        RECT 409.250 191.250 409.750 191.750 ;
        RECT 389.500 190.250 390.000 190.750 ;
        RECT 399.000 190.250 399.500 190.750 ;
        RECT 408.500 190.250 409.000 190.750 ;
        RECT 389.500 189.250 390.000 190.000 ;
        RECT 399.000 189.250 399.500 190.000 ;
        RECT 408.500 189.250 409.000 190.000 ;
        RECT 381.250 188.750 411.250 189.250 ;
        RECT 388.750 187.500 389.250 188.000 ;
        RECT 390.250 187.500 390.750 188.000 ;
        RECT 398.250 187.500 398.750 188.000 ;
        RECT 399.750 187.500 400.250 188.000 ;
        RECT 407.750 187.500 408.250 188.000 ;
        RECT 409.250 187.500 409.750 188.000 ;
        RECT 389.500 186.500 390.000 187.000 ;
        RECT 399.000 186.500 399.500 187.000 ;
        RECT 408.500 186.500 409.000 187.000 ;
        RECT 389.500 185.500 390.000 186.250 ;
        RECT 399.000 185.500 399.500 186.250 ;
        RECT 408.500 185.500 409.000 186.250 ;
        RECT 381.250 185.000 411.250 185.500 ;
        RECT 388.750 183.750 389.250 184.250 ;
        RECT 390.250 183.750 390.750 184.250 ;
        RECT 398.250 183.750 398.750 184.250 ;
        RECT 399.750 183.750 400.250 184.250 ;
        RECT 407.750 183.750 408.250 184.250 ;
        RECT 409.250 183.750 409.750 184.250 ;
        RECT 389.500 182.750 390.000 183.250 ;
        RECT 399.000 182.750 399.500 183.250 ;
        RECT 408.500 182.750 409.000 183.250 ;
        RECT 389.500 181.750 390.000 182.500 ;
        RECT 399.000 181.750 399.500 182.500 ;
        RECT 408.500 181.750 409.000 182.500 ;
        RECT 381.250 181.250 411.250 181.750 ;
        RECT 388.750 180.000 389.250 180.500 ;
        RECT 390.250 180.000 390.750 180.500 ;
        RECT 398.250 180.000 398.750 180.500 ;
        RECT 399.750 180.000 400.250 180.500 ;
        RECT 407.750 180.000 408.250 180.500 ;
        RECT 409.250 180.000 409.750 180.500 ;
        RECT 389.500 179.000 390.000 179.500 ;
        RECT 399.000 179.000 399.500 179.500 ;
        RECT 408.500 179.000 409.000 179.500 ;
        RECT 389.500 178.000 390.000 178.750 ;
        RECT 399.000 178.000 399.500 178.750 ;
        RECT 408.500 178.000 409.000 178.750 ;
        RECT 381.250 177.500 411.250 178.000 ;
        RECT 388.750 176.250 389.250 176.750 ;
        RECT 390.250 176.250 390.750 176.750 ;
        RECT 398.250 176.250 398.750 176.750 ;
        RECT 399.750 176.250 400.250 176.750 ;
        RECT 407.750 176.250 408.250 176.750 ;
        RECT 409.250 176.250 409.750 176.750 ;
        RECT 389.500 175.250 390.000 175.750 ;
        RECT 399.000 175.250 399.500 175.750 ;
        RECT 408.500 175.250 409.000 175.750 ;
        RECT 389.500 174.250 390.000 175.000 ;
        RECT 399.000 174.250 399.500 175.000 ;
        RECT 408.500 174.250 409.000 175.000 ;
        RECT 381.250 173.750 411.250 174.250 ;
        RECT 388.750 172.500 389.250 173.000 ;
        RECT 390.250 172.500 390.750 173.000 ;
        RECT 398.250 172.500 398.750 173.000 ;
        RECT 399.750 172.500 400.250 173.000 ;
        RECT 407.750 172.500 408.250 173.000 ;
        RECT 409.250 172.500 409.750 173.000 ;
        RECT 389.500 171.500 390.000 172.000 ;
        RECT 399.000 171.500 399.500 172.000 ;
        RECT 408.500 171.500 409.000 172.000 ;
        RECT 389.500 170.500 390.000 171.250 ;
        RECT 399.000 170.500 399.500 171.250 ;
        RECT 408.500 170.500 409.000 171.250 ;
        RECT 381.250 170.000 411.250 170.500 ;
        RECT 388.750 168.750 389.250 169.250 ;
        RECT 390.250 168.750 390.750 169.250 ;
        RECT 398.250 168.750 398.750 169.250 ;
        RECT 399.750 168.750 400.250 169.250 ;
        RECT 407.750 168.750 408.250 169.250 ;
        RECT 409.250 168.750 409.750 169.250 ;
        RECT 389.500 167.750 390.000 168.250 ;
        RECT 399.000 167.750 399.500 168.250 ;
        RECT 408.500 167.750 409.000 168.250 ;
        RECT 389.500 166.750 390.000 167.500 ;
        RECT 399.000 166.750 399.500 167.500 ;
        RECT 408.500 166.750 409.000 167.500 ;
        RECT 381.250 166.250 411.250 166.750 ;
        RECT 376.000 152.000 378.000 164.500 ;
        RECT 380.000 157.750 380.500 158.750 ;
        RECT 380.750 153.250 381.750 163.250 ;
        RECT 382.000 157.750 382.500 158.750 ;
        RECT 383.500 157.750 384.000 158.750 ;
        RECT 384.250 153.250 385.250 163.250 ;
        RECT 385.500 157.750 386.000 158.750 ;
        RECT 387.000 157.750 387.500 158.750 ;
        RECT 387.750 153.250 388.750 163.250 ;
        RECT 389.000 157.750 389.500 158.750 ;
        RECT 393.750 156.750 394.250 159.750 ;
        RECT 379.000 109.000 380.000 151.500 ;
        RECT 382.750 150.500 383.750 151.500 ;
        RECT 394.750 150.500 395.750 166.000 ;
        RECT 399.750 156.750 400.250 159.750 ;
        RECT 400.750 150.500 401.750 166.000 ;
        RECT 405.750 156.750 406.250 159.750 ;
        RECT 406.750 150.500 407.750 166.000 ;
        RECT 412.250 163.000 413.250 204.000 ;
        RECT 412.250 156.750 412.750 159.750 ;
        RECT 413.750 156.000 414.250 160.500 ;
        RECT 381.250 149.750 411.250 150.250 ;
        RECT 389.500 149.000 390.000 149.750 ;
        RECT 399.000 149.000 399.500 149.750 ;
        RECT 408.500 149.000 409.000 149.750 ;
        RECT 389.500 148.250 390.000 148.750 ;
        RECT 399.000 148.250 399.500 148.750 ;
        RECT 408.500 148.250 409.000 148.750 ;
        RECT 388.750 147.250 389.250 147.750 ;
        RECT 390.250 147.250 390.750 147.750 ;
        RECT 398.250 147.250 398.750 147.750 ;
        RECT 399.750 147.250 400.250 147.750 ;
        RECT 407.750 147.250 408.250 147.750 ;
        RECT 409.250 147.250 409.750 147.750 ;
        RECT 381.250 146.000 411.250 146.500 ;
        RECT 389.500 145.250 390.000 146.000 ;
        RECT 399.000 145.250 399.500 146.000 ;
        RECT 408.500 145.250 409.000 146.000 ;
        RECT 389.500 144.500 390.000 145.000 ;
        RECT 399.000 144.500 399.500 145.000 ;
        RECT 408.500 144.500 409.000 145.000 ;
        RECT 388.750 143.500 389.250 144.000 ;
        RECT 390.250 143.500 390.750 144.000 ;
        RECT 398.250 143.500 398.750 144.000 ;
        RECT 399.750 143.500 400.250 144.000 ;
        RECT 407.750 143.500 408.250 144.000 ;
        RECT 409.250 143.500 409.750 144.000 ;
        RECT 381.250 142.250 411.250 142.750 ;
        RECT 389.500 141.500 390.000 142.250 ;
        RECT 399.000 141.500 399.500 142.250 ;
        RECT 408.500 141.500 409.000 142.250 ;
        RECT 389.500 140.750 390.000 141.250 ;
        RECT 399.000 140.750 399.500 141.250 ;
        RECT 408.500 140.750 409.000 141.250 ;
        RECT 388.750 139.750 389.250 140.250 ;
        RECT 390.250 139.750 390.750 140.250 ;
        RECT 398.250 139.750 398.750 140.250 ;
        RECT 399.750 139.750 400.250 140.250 ;
        RECT 407.750 139.750 408.250 140.250 ;
        RECT 409.250 139.750 409.750 140.250 ;
        RECT 381.250 138.500 411.250 139.000 ;
        RECT 389.500 137.750 390.000 138.500 ;
        RECT 399.000 137.750 399.500 138.500 ;
        RECT 408.500 137.750 409.000 138.500 ;
        RECT 389.500 137.000 390.000 137.500 ;
        RECT 399.000 137.000 399.500 137.500 ;
        RECT 408.500 137.000 409.000 137.500 ;
        RECT 388.750 136.000 389.250 136.500 ;
        RECT 390.250 136.000 390.750 136.500 ;
        RECT 398.250 136.000 398.750 136.500 ;
        RECT 399.750 136.000 400.250 136.500 ;
        RECT 407.750 136.000 408.250 136.500 ;
        RECT 409.250 136.000 409.750 136.500 ;
        RECT 381.250 134.750 411.250 135.250 ;
        RECT 389.500 134.000 390.000 134.750 ;
        RECT 399.000 134.000 399.500 134.750 ;
        RECT 408.500 134.000 409.000 134.750 ;
        RECT 389.500 133.250 390.000 133.750 ;
        RECT 399.000 133.250 399.500 133.750 ;
        RECT 408.500 133.250 409.000 133.750 ;
        RECT 388.750 132.250 389.250 132.750 ;
        RECT 390.250 132.250 390.750 132.750 ;
        RECT 398.250 132.250 398.750 132.750 ;
        RECT 399.750 132.250 400.250 132.750 ;
        RECT 407.750 132.250 408.250 132.750 ;
        RECT 409.250 132.250 409.750 132.750 ;
        RECT 381.250 131.000 411.250 131.500 ;
        RECT 389.500 130.250 390.000 131.000 ;
        RECT 399.000 130.250 399.500 131.000 ;
        RECT 408.500 130.250 409.000 131.000 ;
        RECT 389.500 129.500 390.000 130.000 ;
        RECT 399.000 129.500 399.500 130.000 ;
        RECT 408.500 129.500 409.000 130.000 ;
        RECT 388.750 128.500 389.250 129.000 ;
        RECT 390.250 128.500 390.750 129.000 ;
        RECT 398.250 128.500 398.750 129.000 ;
        RECT 399.750 128.500 400.250 129.000 ;
        RECT 407.750 128.500 408.250 129.000 ;
        RECT 409.250 128.500 409.750 129.000 ;
        RECT 381.250 127.250 411.250 127.750 ;
        RECT 389.500 126.500 390.000 127.250 ;
        RECT 399.000 126.500 399.500 127.250 ;
        RECT 408.500 126.500 409.000 127.250 ;
        RECT 389.500 125.750 390.000 126.250 ;
        RECT 399.000 125.750 399.500 126.250 ;
        RECT 408.500 125.750 409.000 126.250 ;
        RECT 388.750 124.750 389.250 125.250 ;
        RECT 390.250 124.750 390.750 125.250 ;
        RECT 398.250 124.750 398.750 125.250 ;
        RECT 399.750 124.750 400.250 125.250 ;
        RECT 407.750 124.750 408.250 125.250 ;
        RECT 409.250 124.750 409.750 125.250 ;
        RECT 381.250 123.500 411.250 124.000 ;
        RECT 389.500 122.750 390.000 123.500 ;
        RECT 399.000 122.750 399.500 123.500 ;
        RECT 408.500 122.750 409.000 123.500 ;
        RECT 389.500 122.000 390.000 122.500 ;
        RECT 399.000 122.000 399.500 122.500 ;
        RECT 408.500 122.000 409.000 122.500 ;
        RECT 388.750 121.000 389.250 121.500 ;
        RECT 390.250 121.000 390.750 121.500 ;
        RECT 398.250 121.000 398.750 121.500 ;
        RECT 399.750 121.000 400.250 121.500 ;
        RECT 407.750 121.000 408.250 121.500 ;
        RECT 409.250 121.000 409.750 121.500 ;
        RECT 382.750 109.000 383.750 120.500 ;
        RECT 387.500 109.000 388.500 120.500 ;
        RECT 391.000 109.000 392.000 120.500 ;
        RECT 392.750 119.500 393.250 120.500 ;
        RECT 397.000 109.000 398.000 120.500 ;
        RECT 400.500 109.000 401.500 120.500 ;
        RECT 402.250 119.500 402.750 120.500 ;
        RECT 406.500 109.000 407.500 120.500 ;
        RECT 410.000 109.000 411.000 120.500 ;
        RECT 412.250 109.000 413.250 153.500 ;
        RECT 415.250 104.000 416.500 204.000 ;
        RECT 417.750 156.750 418.250 159.750 ;
        RECT 418.750 152.000 419.750 164.500 ;
      LAYER met3 ;
        RECT 284.500 277.000 306.660 297.400 ;
        RECT 308.000 277.000 330.160 297.400 ;
        RECT 331.500 277.000 353.660 297.400 ;
        RECT 355.000 277.000 377.160 297.400 ;
        RECT 378.500 277.000 400.660 297.400 ;
        RECT 284.500 255.000 306.660 275.400 ;
        RECT 308.000 255.000 330.160 275.400 ;
        RECT 331.500 255.000 353.660 275.400 ;
        RECT 355.000 255.000 377.160 275.400 ;
        RECT 378.500 255.000 400.660 275.400 ;
        RECT 284.500 233.000 306.660 253.400 ;
        RECT 308.000 233.000 330.160 253.400 ;
        RECT 331.500 233.000 353.660 253.400 ;
        RECT 355.000 233.000 377.160 253.400 ;
        RECT 378.500 233.000 400.660 253.400 ;
        RECT 402.000 233.000 424.160 253.400 ;
        RECT 284.500 211.000 306.660 231.400 ;
        RECT 308.000 211.000 330.160 231.400 ;
        RECT 331.500 211.000 353.660 231.400 ;
        RECT 355.000 211.000 377.160 231.400 ;
        RECT 378.500 211.000 400.660 231.400 ;
        RECT 402.000 211.000 424.160 231.400 ;
        RECT 423.000 205.000 427.000 209.000 ;
        RECT 382.750 196.000 383.750 197.000 ;
        RECT 392.750 196.000 393.250 197.000 ;
        RECT 402.250 196.000 402.750 197.000 ;
        RECT 383.250 193.600 387.410 196.000 ;
        RECT 388.750 195.000 389.250 195.500 ;
        RECT 390.250 195.000 390.750 195.500 ;
        RECT 389.500 194.000 391.750 194.500 ;
        RECT 392.750 193.600 396.910 196.000 ;
        RECT 398.250 195.000 398.750 195.500 ;
        RECT 399.750 195.000 400.250 195.500 ;
        RECT 399.000 194.000 401.250 194.500 ;
        RECT 402.250 193.600 406.410 196.000 ;
        RECT 407.750 195.000 408.250 195.500 ;
        RECT 409.250 195.000 409.750 195.500 ;
        RECT 408.500 194.000 410.750 194.500 ;
        RECT 286.500 190.250 325.500 192.250 ;
        RECT 333.750 190.250 350.500 192.250 ;
        RECT 351.500 190.250 353.500 192.250 ;
        RECT 354.500 190.250 358.500 192.250 ;
        RECT 383.250 189.850 387.410 192.250 ;
        RECT 388.750 191.250 389.250 191.750 ;
        RECT 390.250 191.250 390.750 191.750 ;
        RECT 389.500 190.250 391.750 190.750 ;
        RECT 392.750 189.850 396.910 192.250 ;
        RECT 398.250 191.250 398.750 191.750 ;
        RECT 399.750 191.250 400.250 191.750 ;
        RECT 399.000 190.250 401.250 190.750 ;
        RECT 402.250 189.850 406.410 192.250 ;
        RECT 407.750 191.250 408.250 191.750 ;
        RECT 409.250 191.250 409.750 191.750 ;
        RECT 408.500 190.250 410.750 190.750 ;
        RECT 383.250 186.100 387.410 188.500 ;
        RECT 388.750 187.500 389.250 188.000 ;
        RECT 390.250 187.500 390.750 188.000 ;
        RECT 389.500 186.500 391.750 187.000 ;
        RECT 392.750 186.100 396.910 188.500 ;
        RECT 398.250 187.500 398.750 188.000 ;
        RECT 399.750 187.500 400.250 188.000 ;
        RECT 399.000 186.500 401.250 187.000 ;
        RECT 402.250 186.100 406.410 188.500 ;
        RECT 407.750 187.500 408.250 188.000 ;
        RECT 409.250 187.500 409.750 188.000 ;
        RECT 408.500 186.500 410.750 187.000 ;
        RECT 285.500 183.100 289.500 183.500 ;
        RECT 296.765 183.100 297.095 183.115 ;
        RECT 285.500 182.800 297.095 183.100 ;
        RECT 285.500 182.500 289.500 182.800 ;
        RECT 296.765 182.785 297.095 182.800 ;
        RECT 300.460 183.100 300.790 183.115 ;
        RECT 319.250 183.100 360.000 183.500 ;
        RECT 300.460 182.800 360.000 183.100 ;
        RECT 300.460 182.785 300.790 182.800 ;
        RECT 319.250 182.500 360.000 182.800 ;
        RECT 383.250 182.350 387.410 184.750 ;
        RECT 388.750 183.750 389.250 184.250 ;
        RECT 390.250 183.750 390.750 184.250 ;
        RECT 389.500 182.750 391.750 183.250 ;
        RECT 392.750 182.350 396.910 184.750 ;
        RECT 398.250 183.750 398.750 184.250 ;
        RECT 399.750 183.750 400.250 184.250 ;
        RECT 399.000 182.750 401.250 183.250 ;
        RECT 402.250 182.350 406.410 184.750 ;
        RECT 407.750 183.750 408.250 184.250 ;
        RECT 409.250 183.750 409.750 184.250 ;
        RECT 408.500 182.750 410.750 183.250 ;
        RECT 285.500 181.600 289.500 182.000 ;
        RECT 296.305 181.600 296.635 181.615 ;
        RECT 285.500 181.300 296.635 181.600 ;
        RECT 285.500 181.000 289.500 181.300 ;
        RECT 296.305 181.285 296.635 181.300 ;
        RECT 297.685 181.600 298.015 181.615 ;
        RECT 319.250 181.600 361.000 182.000 ;
        RECT 297.685 181.300 361.000 181.600 ;
        RECT 297.685 181.285 298.015 181.300 ;
        RECT 319.250 181.000 361.000 181.300 ;
        RECT 285.500 180.100 289.500 180.500 ;
        RECT 311.850 180.475 313.430 180.805 ;
        RECT 299.985 180.100 300.315 180.115 ;
        RECT 285.500 179.800 300.315 180.100 ;
        RECT 285.500 179.500 289.500 179.800 ;
        RECT 299.985 179.785 300.315 179.800 ;
        RECT 300.935 180.100 301.265 180.115 ;
        RECT 319.250 180.100 362.000 180.500 ;
        RECT 300.935 179.800 362.000 180.100 ;
        RECT 300.935 179.785 301.265 179.800 ;
        RECT 319.250 179.500 362.000 179.800 ;
        RECT 285.500 178.600 289.500 179.000 ;
        RECT 297.225 178.600 297.555 178.615 ;
        RECT 285.500 178.300 297.555 178.600 ;
        RECT 285.500 178.000 289.500 178.300 ;
        RECT 297.225 178.285 297.555 178.300 ;
        RECT 301.410 178.600 301.740 178.615 ;
        RECT 319.250 178.600 363.000 179.000 ;
        RECT 383.250 178.600 387.410 181.000 ;
        RECT 388.750 180.000 389.250 180.500 ;
        RECT 390.250 180.000 390.750 180.500 ;
        RECT 389.500 179.000 391.750 179.500 ;
        RECT 392.750 178.600 396.910 181.000 ;
        RECT 398.250 180.000 398.750 180.500 ;
        RECT 399.750 180.000 400.250 180.500 ;
        RECT 399.000 179.000 401.250 179.500 ;
        RECT 402.250 178.600 406.410 181.000 ;
        RECT 407.750 180.000 408.250 180.500 ;
        RECT 409.250 180.000 409.750 180.500 ;
        RECT 408.500 179.000 410.750 179.500 ;
        RECT 301.410 178.300 363.000 178.600 ;
        RECT 301.410 178.285 301.740 178.300 ;
        RECT 319.250 178.000 363.000 178.300 ;
        RECT 313.785 177.100 314.115 177.115 ;
        RECT 319.250 177.100 364.000 177.500 ;
        RECT 313.785 176.800 364.000 177.100 ;
        RECT 313.785 176.785 314.115 176.800 ;
        RECT 319.250 176.500 364.000 176.800 ;
        RECT 314.245 175.600 314.575 175.615 ;
        RECT 319.250 175.600 365.000 176.000 ;
        RECT 314.245 175.300 365.000 175.600 ;
        RECT 314.245 175.285 314.575 175.300 ;
        RECT 319.250 175.000 365.000 175.300 ;
        RECT 383.250 174.850 387.410 177.250 ;
        RECT 388.750 176.250 389.250 176.750 ;
        RECT 390.250 176.250 390.750 176.750 ;
        RECT 389.500 175.250 391.750 175.750 ;
        RECT 392.750 174.850 396.910 177.250 ;
        RECT 398.250 176.250 398.750 176.750 ;
        RECT 399.750 176.250 400.250 176.750 ;
        RECT 399.000 175.250 401.250 175.750 ;
        RECT 402.250 174.850 406.410 177.250 ;
        RECT 407.750 176.250 408.250 176.750 ;
        RECT 409.250 176.250 409.750 176.750 ;
        RECT 408.500 175.250 410.750 175.750 ;
        RECT 314.705 174.100 315.035 174.115 ;
        RECT 319.250 174.100 366.000 174.500 ;
        RECT 314.705 173.800 366.000 174.100 ;
        RECT 314.705 173.785 315.035 173.800 ;
        RECT 319.250 173.500 366.000 173.800 ;
        RECT 313.325 172.600 313.655 172.615 ;
        RECT 319.250 172.600 367.000 173.000 ;
        RECT 313.325 172.300 367.000 172.600 ;
        RECT 313.325 172.285 313.655 172.300 ;
        RECT 319.250 172.000 367.000 172.300 ;
        RECT 317.005 171.100 317.335 171.115 ;
        RECT 319.250 171.100 368.000 171.500 ;
        RECT 383.250 171.100 387.410 173.500 ;
        RECT 388.750 172.500 389.250 173.000 ;
        RECT 390.250 172.500 390.750 173.000 ;
        RECT 389.500 171.500 391.750 172.000 ;
        RECT 392.750 171.100 396.910 173.500 ;
        RECT 398.250 172.500 398.750 173.000 ;
        RECT 399.750 172.500 400.250 173.000 ;
        RECT 399.000 171.500 401.250 172.000 ;
        RECT 402.250 171.100 406.410 173.500 ;
        RECT 407.750 172.500 408.250 173.000 ;
        RECT 409.250 172.500 409.750 173.000 ;
        RECT 408.500 171.500 410.750 172.000 ;
        RECT 317.005 170.800 368.000 171.100 ;
        RECT 317.005 170.785 317.335 170.800 ;
        RECT 319.250 170.500 368.000 170.800 ;
        RECT 312.865 169.600 313.195 169.615 ;
        RECT 319.250 169.600 369.000 170.000 ;
        RECT 312.865 169.300 369.000 169.600 ;
        RECT 312.865 169.285 313.195 169.300 ;
        RECT 319.250 169.000 369.000 169.300 ;
        RECT 295.845 168.100 296.175 168.115 ;
        RECT 319.250 168.100 370.000 168.500 ;
        RECT 295.845 167.800 370.000 168.100 ;
        RECT 295.845 167.785 296.175 167.800 ;
        RECT 319.250 167.500 370.000 167.800 ;
        RECT 383.250 167.350 387.410 169.750 ;
        RECT 388.750 168.750 389.250 169.250 ;
        RECT 390.250 168.750 390.750 169.250 ;
        RECT 389.500 167.750 391.750 168.250 ;
        RECT 392.750 167.350 396.910 169.750 ;
        RECT 398.250 168.750 398.750 169.250 ;
        RECT 399.750 168.750 400.250 169.250 ;
        RECT 399.000 167.750 401.250 168.250 ;
        RECT 402.250 167.350 406.410 169.750 ;
        RECT 407.750 168.750 408.250 169.250 ;
        RECT 409.250 168.750 409.750 169.250 ;
        RECT 408.500 167.750 410.750 168.250 ;
        RECT 297.685 166.600 298.015 166.615 ;
        RECT 319.250 166.600 371.000 167.000 ;
        RECT 297.685 166.300 371.000 166.600 ;
        RECT 297.685 166.285 298.015 166.300 ;
        RECT 319.250 166.000 371.000 166.300 ;
        RECT 295.385 165.100 295.715 165.115 ;
        RECT 319.250 165.100 372.000 165.500 ;
        RECT 295.385 164.800 372.000 165.100 ;
        RECT 391.250 165.000 395.750 166.000 ;
        RECT 400.750 165.000 401.750 166.000 ;
        RECT 406.750 165.000 411.250 166.000 ;
        RECT 295.385 164.785 295.715 164.800 ;
        RECT 319.250 164.500 372.000 164.800 ;
        RECT 300.445 163.700 300.775 163.715 ;
        RECT 319.250 163.700 373.000 164.000 ;
        RECT 376.000 163.750 419.750 164.500 ;
        RECT 300.445 163.400 373.000 163.700 ;
        RECT 300.445 163.385 300.775 163.400 ;
        RECT 319.250 163.000 373.000 163.400 ;
        RECT 381.250 162.750 395.250 163.250 ;
        RECT 299.525 162.100 299.855 162.115 ;
        RECT 319.250 162.100 374.000 162.500 ;
        RECT 299.525 161.800 374.000 162.100 ;
        RECT 299.525 161.785 299.855 161.800 ;
        RECT 319.250 161.500 374.000 161.800 ;
        RECT 384.750 161.750 401.250 162.250 ;
        RECT 294.465 160.600 294.795 160.615 ;
        RECT 319.250 160.600 375.000 161.000 ;
        RECT 388.250 160.750 407.250 161.250 ;
        RECT 294.465 160.300 375.000 160.600 ;
        RECT 294.465 160.285 294.795 160.300 ;
        RECT 319.250 160.000 375.000 160.300 ;
        RECT 393.750 159.250 407.250 159.750 ;
        RECT 299.250 156.000 301.250 158.000 ;
        RECT 356.500 157.500 376.000 159.000 ;
        RECT 377.500 157.500 389.500 159.000 ;
        RECT 419.250 158.750 422.500 159.250 ;
        RECT 395.250 158.000 400.250 158.500 ;
        RECT 401.250 158.000 406.250 158.500 ;
        RECT 407.250 158.000 412.750 158.500 ;
        RECT 413.750 158.000 418.250 158.500 ;
        RECT 418.750 157.750 422.500 158.750 ;
        RECT 419.250 157.250 422.500 157.750 ;
        RECT 393.750 156.750 407.250 157.250 ;
        RECT 388.250 155.250 407.250 155.750 ;
        RECT 384.750 154.250 401.250 154.750 ;
        RECT 381.250 153.250 395.250 153.750 ;
        RECT 376.000 152.000 419.750 152.750 ;
        RECT 382.750 150.500 383.750 151.500 ;
        RECT 391.250 150.500 395.750 151.500 ;
        RECT 400.750 150.500 401.750 151.500 ;
        RECT 406.750 150.500 411.250 151.500 ;
        RECT 285.500 149.500 339.000 150.500 ;
        RECT 285.500 148.000 326.000 149.000 ;
        RECT 285.500 146.500 318.500 147.500 ;
        RECT 383.250 146.750 387.410 149.150 ;
        RECT 389.500 148.250 391.750 148.750 ;
        RECT 388.750 147.250 389.250 147.750 ;
        RECT 390.250 147.250 390.750 147.750 ;
        RECT 392.750 146.750 396.910 149.150 ;
        RECT 399.000 148.250 401.250 148.750 ;
        RECT 398.250 147.250 398.750 147.750 ;
        RECT 399.750 147.250 400.250 147.750 ;
        RECT 402.250 146.750 406.410 149.150 ;
        RECT 408.500 148.250 410.750 148.750 ;
        RECT 407.750 147.250 408.250 147.750 ;
        RECT 409.250 147.250 409.750 147.750 ;
        RECT 285.500 145.000 331.500 146.000 ;
        RECT 383.250 143.000 387.410 145.400 ;
        RECT 389.500 144.500 391.750 145.000 ;
        RECT 388.750 143.500 389.250 144.000 ;
        RECT 390.250 143.500 390.750 144.000 ;
        RECT 392.750 143.000 396.910 145.400 ;
        RECT 399.000 144.500 401.250 145.000 ;
        RECT 398.250 143.500 398.750 144.000 ;
        RECT 399.750 143.500 400.250 144.000 ;
        RECT 402.250 143.000 406.410 145.400 ;
        RECT 408.500 144.500 410.750 145.000 ;
        RECT 407.750 143.500 408.250 144.000 ;
        RECT 409.250 143.500 409.750 144.000 ;
        RECT 303.500 138.750 304.000 139.250 ;
        RECT 304.500 137.000 309.750 141.400 ;
        RECT 311.000 137.000 316.250 141.400 ;
        RECT 325.000 138.500 326.000 139.500 ;
        RECT 338.000 138.500 339.000 139.500 ;
        RECT 383.250 139.250 387.410 141.650 ;
        RECT 389.500 140.750 391.750 141.250 ;
        RECT 388.750 139.750 389.250 140.250 ;
        RECT 390.250 139.750 390.750 140.250 ;
        RECT 392.750 139.250 396.910 141.650 ;
        RECT 399.000 140.750 401.250 141.250 ;
        RECT 398.250 139.750 398.750 140.250 ;
        RECT 399.750 139.750 400.250 140.250 ;
        RECT 402.250 139.250 406.410 141.650 ;
        RECT 408.500 140.750 410.750 141.250 ;
        RECT 407.750 139.750 408.250 140.250 ;
        RECT 409.250 139.750 409.750 140.250 ;
        RECT 383.250 135.500 387.410 137.900 ;
        RECT 389.500 137.000 391.750 137.500 ;
        RECT 388.750 136.000 389.250 136.500 ;
        RECT 390.250 136.000 390.750 136.500 ;
        RECT 392.750 135.500 396.910 137.900 ;
        RECT 399.000 137.000 401.250 137.500 ;
        RECT 398.250 136.000 398.750 136.500 ;
        RECT 399.750 136.000 400.250 136.500 ;
        RECT 402.250 135.500 406.410 137.900 ;
        RECT 408.500 137.000 410.750 137.500 ;
        RECT 407.750 136.000 408.250 136.500 ;
        RECT 409.250 136.000 409.750 136.500 ;
        RECT 303.500 131.750 304.000 132.250 ;
        RECT 304.500 130.000 309.750 134.400 ;
        RECT 311.750 131.750 313.000 132.250 ;
        RECT 317.500 131.500 318.500 132.500 ;
        RECT 330.500 131.500 331.500 132.500 ;
        RECT 383.250 131.750 387.410 134.150 ;
        RECT 389.500 133.250 391.750 133.750 ;
        RECT 388.750 132.250 389.250 132.750 ;
        RECT 390.250 132.250 390.750 132.750 ;
        RECT 392.750 131.750 396.910 134.150 ;
        RECT 399.000 133.250 401.250 133.750 ;
        RECT 398.250 132.250 398.750 132.750 ;
        RECT 399.750 132.250 400.250 132.750 ;
        RECT 402.250 131.750 406.410 134.150 ;
        RECT 408.500 133.250 410.750 133.750 ;
        RECT 407.750 132.250 408.250 132.750 ;
        RECT 409.250 132.250 409.750 132.750 ;
        RECT 383.250 128.000 387.410 130.400 ;
        RECT 389.500 129.500 391.750 130.000 ;
        RECT 388.750 128.500 389.250 129.000 ;
        RECT 390.250 128.500 390.750 129.000 ;
        RECT 392.750 128.000 396.910 130.400 ;
        RECT 399.000 129.500 401.250 130.000 ;
        RECT 398.250 128.500 398.750 129.000 ;
        RECT 399.750 128.500 400.250 129.000 ;
        RECT 402.250 128.000 406.410 130.400 ;
        RECT 408.500 129.500 410.750 130.000 ;
        RECT 407.750 128.500 408.250 129.000 ;
        RECT 409.250 128.500 409.750 129.000 ;
        RECT 383.250 124.250 387.410 126.650 ;
        RECT 389.500 125.750 391.750 126.250 ;
        RECT 388.750 124.750 389.250 125.250 ;
        RECT 390.250 124.750 390.750 125.250 ;
        RECT 392.750 124.250 396.910 126.650 ;
        RECT 399.000 125.750 401.250 126.250 ;
        RECT 398.250 124.750 398.750 125.250 ;
        RECT 399.750 124.750 400.250 125.250 ;
        RECT 402.250 124.250 406.410 126.650 ;
        RECT 408.500 125.750 410.750 126.250 ;
        RECT 407.750 124.750 408.250 125.250 ;
        RECT 409.250 124.750 409.750 125.250 ;
        RECT 285.500 119.750 344.000 120.750 ;
        RECT 383.250 120.500 387.410 122.900 ;
        RECT 389.500 122.000 391.750 122.500 ;
        RECT 388.750 121.000 389.250 121.500 ;
        RECT 390.250 121.000 390.750 121.500 ;
        RECT 392.750 120.500 396.910 122.900 ;
        RECT 399.000 122.000 401.250 122.500 ;
        RECT 398.250 121.000 398.750 121.500 ;
        RECT 399.750 121.000 400.250 121.500 ;
        RECT 402.250 120.500 406.410 122.900 ;
        RECT 408.500 122.000 410.750 122.500 ;
        RECT 407.750 121.000 408.250 121.500 ;
        RECT 409.250 121.000 409.750 121.500 ;
        RECT 382.750 119.500 383.750 120.500 ;
        RECT 392.750 119.500 393.250 120.500 ;
        RECT 402.250 119.500 402.750 120.500 ;
        RECT 285.500 117.750 338.000 118.750 ;
        RECT 299.250 115.750 308.250 116.750 ;
      LAYER met4 ;
        RECT 305.500 298.000 425.000 300.000 ;
        RECT 293.500 297.005 295.500 297.500 ;
        RECT 284.895 277.395 304.505 297.005 ;
        RECT 293.500 275.005 295.500 277.395 ;
        RECT 284.895 255.395 304.505 275.005 ;
        RECT 293.500 253.005 295.500 255.395 ;
        RECT 284.895 233.395 304.505 253.005 ;
        RECT 293.500 231.005 295.500 233.395 ;
        RECT 284.895 211.395 304.505 231.005 ;
        RECT 293.500 210.500 295.500 211.395 ;
        RECT 305.500 211.000 307.500 298.000 ;
        RECT 317.000 297.005 319.000 297.500 ;
        RECT 308.395 277.395 328.005 297.005 ;
        RECT 317.000 275.005 319.000 277.395 ;
        RECT 308.395 255.395 328.005 275.005 ;
        RECT 317.000 253.005 319.000 255.395 ;
        RECT 308.395 233.395 328.005 253.005 ;
        RECT 317.000 231.005 319.000 233.395 ;
        RECT 308.395 211.395 328.005 231.005 ;
        RECT 317.000 210.500 319.000 211.395 ;
        RECT 329.000 211.000 331.000 298.000 ;
        RECT 340.500 297.005 342.500 297.500 ;
        RECT 331.895 277.395 351.505 297.005 ;
        RECT 340.500 275.005 342.500 277.395 ;
        RECT 331.895 255.395 351.505 275.005 ;
        RECT 340.500 253.005 342.500 255.395 ;
        RECT 331.895 233.395 351.505 253.005 ;
        RECT 340.500 231.005 342.500 233.395 ;
        RECT 331.895 211.395 351.505 231.005 ;
        RECT 340.500 210.500 342.500 211.395 ;
        RECT 352.500 211.000 354.500 298.000 ;
        RECT 364.000 297.005 366.000 297.500 ;
        RECT 355.395 277.395 375.005 297.005 ;
        RECT 364.000 275.005 366.000 277.395 ;
        RECT 355.395 255.395 375.005 275.005 ;
        RECT 364.000 253.005 366.000 255.395 ;
        RECT 355.395 233.395 375.005 253.005 ;
        RECT 364.000 231.005 366.000 233.395 ;
        RECT 355.395 211.395 375.005 231.005 ;
        RECT 364.000 210.500 366.000 211.395 ;
        RECT 376.000 211.000 378.000 298.000 ;
        RECT 387.500 297.005 389.500 297.500 ;
        RECT 378.895 277.395 398.505 297.005 ;
        RECT 387.500 275.005 389.500 277.395 ;
        RECT 378.895 255.395 398.505 275.005 ;
        RECT 387.500 253.005 389.500 255.395 ;
        RECT 378.895 233.395 398.505 253.005 ;
        RECT 387.500 231.005 389.500 233.395 ;
        RECT 378.895 211.395 398.505 231.005 ;
        RECT 387.500 210.500 389.500 211.395 ;
        RECT 399.500 211.000 401.500 298.000 ;
        RECT 411.000 253.005 413.000 253.500 ;
        RECT 402.395 233.395 422.005 253.005 ;
        RECT 411.000 231.005 413.000 233.395 ;
        RECT 402.395 211.395 422.005 231.005 ;
        RECT 293.500 208.500 389.500 210.500 ;
        RECT 351.250 189.500 353.750 208.500 ;
        RECT 411.000 208.000 413.000 211.395 ;
        RECT 356.500 206.000 413.000 208.000 ;
        RECT 423.000 209.000 425.000 298.000 ;
        RECT 299.250 115.750 301.250 158.000 ;
        RECT 356.500 157.500 358.500 206.000 ;
        RECT 423.000 205.000 427.000 209.000 ;
        RECT 305.745 139.250 309.355 141.005 ;
        RECT 303.500 138.750 309.355 139.250 ;
        RECT 305.745 137.395 309.355 138.750 ;
        RECT 312.245 137.395 315.855 141.005 ;
        RECT 305.745 132.250 309.355 134.005 ;
        RECT 303.500 131.750 309.355 132.250 ;
        RECT 312.500 131.750 313.000 137.395 ;
        RECT 305.745 130.395 309.355 131.750 ;
        RECT 317.500 131.500 318.500 147.500 ;
        RECT 325.000 138.500 326.000 149.000 ;
        RECT 330.500 131.500 331.500 146.000 ;
        RECT 338.000 138.500 339.000 150.500 ;
        RECT 382.750 119.500 383.750 197.000 ;
        RECT 385.405 195.500 387.015 195.605 ;
        RECT 385.405 195.000 390.750 195.500 ;
        RECT 385.405 193.995 387.015 195.000 ;
        RECT 385.405 191.750 387.015 191.855 ;
        RECT 385.405 191.250 390.750 191.750 ;
        RECT 385.405 190.245 387.015 191.250 ;
        RECT 385.405 188.000 387.015 188.105 ;
        RECT 385.405 187.500 390.750 188.000 ;
        RECT 385.405 186.495 387.015 187.500 ;
        RECT 385.405 184.250 387.015 184.355 ;
        RECT 385.405 183.750 390.750 184.250 ;
        RECT 385.405 182.745 387.015 183.750 ;
        RECT 385.405 180.500 387.015 180.605 ;
        RECT 385.405 180.000 390.750 180.500 ;
        RECT 385.405 178.995 387.015 180.000 ;
        RECT 385.405 176.750 387.015 176.855 ;
        RECT 385.405 176.250 390.750 176.750 ;
        RECT 385.405 175.245 387.015 176.250 ;
        RECT 385.405 173.000 387.015 173.105 ;
        RECT 385.405 172.500 390.750 173.000 ;
        RECT 385.405 171.495 387.015 172.500 ;
        RECT 385.405 169.250 387.015 169.355 ;
        RECT 385.405 168.750 390.750 169.250 ;
        RECT 385.405 167.745 387.015 168.750 ;
        RECT 391.250 165.000 392.250 194.500 ;
        RECT 392.750 167.250 393.250 197.000 ;
        RECT 394.905 195.500 396.515 195.605 ;
        RECT 394.905 195.000 400.250 195.500 ;
        RECT 394.905 193.995 396.515 195.000 ;
        RECT 394.905 191.750 396.515 191.855 ;
        RECT 394.905 191.250 400.250 191.750 ;
        RECT 394.905 190.245 396.515 191.250 ;
        RECT 394.905 188.000 396.515 188.105 ;
        RECT 394.905 187.500 400.250 188.000 ;
        RECT 394.905 186.495 396.515 187.500 ;
        RECT 394.905 184.250 396.515 184.355 ;
        RECT 394.905 183.750 400.250 184.250 ;
        RECT 394.905 182.745 396.515 183.750 ;
        RECT 394.905 180.500 396.515 180.605 ;
        RECT 394.905 180.000 400.250 180.500 ;
        RECT 394.905 178.995 396.515 180.000 ;
        RECT 394.905 176.750 396.515 176.855 ;
        RECT 394.905 176.250 400.250 176.750 ;
        RECT 394.905 175.245 396.515 176.250 ;
        RECT 394.905 173.000 396.515 173.105 ;
        RECT 394.905 172.500 400.250 173.000 ;
        RECT 394.905 171.495 396.515 172.500 ;
        RECT 394.905 169.250 396.515 169.355 ;
        RECT 394.905 168.750 400.250 169.250 ;
        RECT 394.905 167.745 396.515 168.750 ;
        RECT 400.750 165.000 401.750 194.500 ;
        RECT 402.250 167.250 402.750 197.000 ;
        RECT 404.405 195.500 406.015 195.605 ;
        RECT 404.405 195.000 409.750 195.500 ;
        RECT 404.405 193.995 406.015 195.000 ;
        RECT 404.405 191.750 406.015 191.855 ;
        RECT 404.405 191.250 409.750 191.750 ;
        RECT 404.405 190.245 406.015 191.250 ;
        RECT 404.405 188.000 406.015 188.105 ;
        RECT 404.405 187.500 409.750 188.000 ;
        RECT 404.405 186.495 406.015 187.500 ;
        RECT 404.405 184.250 406.015 184.355 ;
        RECT 404.405 183.750 409.750 184.250 ;
        RECT 404.405 182.745 406.015 183.750 ;
        RECT 404.405 180.500 406.015 180.605 ;
        RECT 404.405 180.000 409.750 180.500 ;
        RECT 404.405 178.995 406.015 180.000 ;
        RECT 404.405 176.750 406.015 176.855 ;
        RECT 404.405 176.250 409.750 176.750 ;
        RECT 404.405 175.245 406.015 176.250 ;
        RECT 404.405 173.000 406.015 173.105 ;
        RECT 404.405 172.500 409.750 173.000 ;
        RECT 404.405 171.495 406.015 172.500 ;
        RECT 404.405 169.250 406.015 169.355 ;
        RECT 404.405 168.750 409.750 169.250 ;
        RECT 404.405 167.745 406.015 168.750 ;
        RECT 410.250 165.000 411.250 194.500 ;
        RECT 385.405 147.750 387.015 148.755 ;
        RECT 385.405 147.250 390.750 147.750 ;
        RECT 385.405 147.145 387.015 147.250 ;
        RECT 385.405 144.000 387.015 145.005 ;
        RECT 385.405 143.500 390.750 144.000 ;
        RECT 385.405 143.395 387.015 143.500 ;
        RECT 385.405 140.250 387.015 141.255 ;
        RECT 385.405 139.750 390.750 140.250 ;
        RECT 385.405 139.645 387.015 139.750 ;
        RECT 385.405 136.500 387.015 137.505 ;
        RECT 385.405 136.000 390.750 136.500 ;
        RECT 385.405 135.895 387.015 136.000 ;
        RECT 385.405 132.750 387.015 133.755 ;
        RECT 385.405 132.250 390.750 132.750 ;
        RECT 385.405 132.145 387.015 132.250 ;
        RECT 385.405 129.000 387.015 130.005 ;
        RECT 385.405 128.500 390.750 129.000 ;
        RECT 385.405 128.395 387.015 128.500 ;
        RECT 385.405 125.250 387.015 126.255 ;
        RECT 385.405 124.750 390.750 125.250 ;
        RECT 385.405 124.645 387.015 124.750 ;
        RECT 385.405 121.500 387.015 122.505 ;
        RECT 391.250 122.000 392.250 151.500 ;
        RECT 385.405 121.000 390.750 121.500 ;
        RECT 385.405 120.895 387.015 121.000 ;
        RECT 392.750 119.500 393.250 149.250 ;
        RECT 394.905 147.750 396.515 148.755 ;
        RECT 394.905 147.250 400.250 147.750 ;
        RECT 394.905 147.145 396.515 147.250 ;
        RECT 394.905 144.000 396.515 145.005 ;
        RECT 394.905 143.500 400.250 144.000 ;
        RECT 394.905 143.395 396.515 143.500 ;
        RECT 394.905 140.250 396.515 141.255 ;
        RECT 394.905 139.750 400.250 140.250 ;
        RECT 394.905 139.645 396.515 139.750 ;
        RECT 394.905 136.500 396.515 137.505 ;
        RECT 394.905 136.000 400.250 136.500 ;
        RECT 394.905 135.895 396.515 136.000 ;
        RECT 394.905 132.750 396.515 133.755 ;
        RECT 394.905 132.250 400.250 132.750 ;
        RECT 394.905 132.145 396.515 132.250 ;
        RECT 394.905 129.000 396.515 130.005 ;
        RECT 394.905 128.500 400.250 129.000 ;
        RECT 394.905 128.395 396.515 128.500 ;
        RECT 394.905 125.250 396.515 126.255 ;
        RECT 394.905 124.750 400.250 125.250 ;
        RECT 394.905 124.645 396.515 124.750 ;
        RECT 394.905 121.500 396.515 122.505 ;
        RECT 400.750 122.000 401.750 151.500 ;
        RECT 394.905 121.000 400.250 121.500 ;
        RECT 394.905 120.895 396.515 121.000 ;
        RECT 402.250 119.500 402.750 149.250 ;
        RECT 404.405 147.750 406.015 148.755 ;
        RECT 404.405 147.250 409.750 147.750 ;
        RECT 404.405 147.145 406.015 147.250 ;
        RECT 404.405 144.000 406.015 145.005 ;
        RECT 404.405 143.500 409.750 144.000 ;
        RECT 404.405 143.395 406.015 143.500 ;
        RECT 404.405 140.250 406.015 141.255 ;
        RECT 404.405 139.750 409.750 140.250 ;
        RECT 404.405 139.645 406.015 139.750 ;
        RECT 404.405 136.500 406.015 137.505 ;
        RECT 404.405 136.000 409.750 136.500 ;
        RECT 404.405 135.895 406.015 136.000 ;
        RECT 404.405 132.750 406.015 133.755 ;
        RECT 404.405 132.250 409.750 132.750 ;
        RECT 404.405 132.145 406.015 132.250 ;
        RECT 404.405 129.000 406.015 130.005 ;
        RECT 404.405 128.500 409.750 129.000 ;
        RECT 404.405 128.395 406.015 128.500 ;
        RECT 404.405 125.250 406.015 126.255 ;
        RECT 404.405 124.750 409.750 125.250 ;
        RECT 404.405 124.645 406.015 124.750 ;
        RECT 404.405 121.500 406.015 122.505 ;
        RECT 410.250 122.000 411.250 151.500 ;
        RECT 404.405 121.000 409.750 121.500 ;
        RECT 404.405 120.895 406.015 121.000 ;
  END
END tl_synth_v4
END LIBRARY

